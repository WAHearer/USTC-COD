
`timescale 1ns/1ps
module mem_bram #(
    parameter ADDR_WIDTH = 10,		//地址宽度
    parameter DATA_WIDTH = 128		//数据宽度
)(
    input                   clk,   // Clock
    input [ADDR_WIDTH-1:0]  raddr,  // Address
    input [ADDR_WIDTH-1:0]  waddr,  // Address
    input [DATA_WIDTH-1:0]  din,   // Data Input
    input                   we,    // Write Enable
    output [DATA_WIDTH-1:0] dout   // Data Output
); 
    reg [ADDR_WIDTH-1:0] addr_r;  // Address Register
    reg [DATA_WIDTH-1:0] ram [0:(1 << ADDR_WIDTH)-1];
    integer i;
    initial begin
        ram[0][31:0] = 32'd1241483398;
        ram[0][63:32] = 32'd1830337710;
        ram[0][95:64] = 32'd2722018698;
        ram[0][127:96] = 32'd3665711875;
        ram[1][31:0] = 32'd340910773;
        ram[1][63:32] = 32'd426215752;
        ram[1][95:64] = 32'd805363560;
        ram[1][127:96] = 32'd721822125;
        ram[2][31:0] = 32'd4176320574;
        ram[2][63:32] = 32'd3430358658;
        ram[2][95:64] = 32'd3074773431;
        ram[2][127:96] = 32'd1390075433;
        ram[3][31:0] = 32'd1442523325;
        ram[3][63:32] = 32'd2440374455;
        ram[3][95:64] = 32'd1328303385;
        ram[3][127:96] = 32'd2428622533;
        ram[4][31:0] = 32'd38352283;
        ram[4][63:32] = 32'd3107376114;
        ram[4][95:64] = 32'd677422689;
        ram[4][127:96] = 32'd3066389384;
        ram[5][31:0] = 32'd2974051818;
        ram[5][63:32] = 32'd513590475;
        ram[5][95:64] = 32'd3991520861;
        ram[5][127:96] = 32'd860970747;
        ram[6][31:0] = 32'd759408867;
        ram[6][63:32] = 32'd2632895408;
        ram[6][95:64] = 32'd3295931461;
        ram[6][127:96] = 32'd1081001156;
        ram[7][31:0] = 32'd1285008039;
        ram[7][63:32] = 32'd943496892;
        ram[7][95:64] = 32'd393122722;
        ram[7][127:96] = 32'd3195599876;
        ram[8][31:0] = 32'd4281965901;
        ram[8][63:32] = 32'd3213587532;
        ram[8][95:64] = 32'd3363095958;
        ram[8][127:96] = 32'd1763527796;
        ram[9][31:0] = 32'd2630607988;
        ram[9][63:32] = 32'd2923110415;
        ram[9][95:64] = 32'd849503955;
        ram[9][127:96] = 32'd2019161959;
        ram[10][31:0] = 32'd2719542166;
        ram[10][63:32] = 32'd1144135439;
        ram[10][95:64] = 32'd3158623633;
        ram[10][127:96] = 32'd2969307118;
        ram[11][31:0] = 32'd3264450694;
        ram[11][63:32] = 32'd3609312874;
        ram[11][95:64] = 32'd1283596394;
        ram[11][127:96] = 32'd1960792394;
        ram[12][31:0] = 32'd3555854734;
        ram[12][63:32] = 32'd3795521150;
        ram[12][95:64] = 32'd3517050998;
        ram[12][127:96] = 32'd3196449230;
        ram[13][31:0] = 32'd1670309798;
        ram[13][63:32] = 32'd150061981;
        ram[13][95:64] = 32'd586437743;
        ram[13][127:96] = 32'd1399484111;
        ram[14][31:0] = 32'd4032767092;
        ram[14][63:32] = 32'd3015078990;
        ram[14][95:64] = 32'd2630100688;
        ram[14][127:96] = 32'd3954950459;
        ram[15][31:0] = 32'd132987420;
        ram[15][63:32] = 32'd2025170720;
        ram[15][95:64] = 32'd304754323;
        ram[15][127:96] = 32'd1646915880;
        ram[16][31:0] = 32'd2718552178;
        ram[16][63:32] = 32'd1845517365;
        ram[16][95:64] = 32'd2814571527;
        ram[16][127:96] = 32'd1049063200;
        ram[17][31:0] = 32'd2448672930;
        ram[17][63:32] = 32'd1109676571;
        ram[17][95:64] = 32'd2049921272;
        ram[17][127:96] = 32'd2763155768;
        ram[18][31:0] = 32'd46563330;
        ram[18][63:32] = 32'd404406686;
        ram[18][95:64] = 32'd3957199885;
        ram[18][127:96] = 32'd869866033;
        ram[19][31:0] = 32'd1934095929;
        ram[19][63:32] = 32'd2876543838;
        ram[19][95:64] = 32'd3671955214;
        ram[19][127:96] = 32'd238733017;
        ram[20][31:0] = 32'd2907114715;
        ram[20][63:32] = 32'd1759133022;
        ram[20][95:64] = 32'd2394041630;
        ram[20][127:96] = 32'd21120565;
        ram[21][31:0] = 32'd655204540;
        ram[21][63:32] = 32'd4049262913;
        ram[21][95:64] = 32'd88473128;
        ram[21][127:96] = 32'd1351154336;
        ram[22][31:0] = 32'd2644571144;
        ram[22][63:32] = 32'd227902140;
        ram[22][95:64] = 32'd222554208;
        ram[22][127:96] = 32'd2419969866;
        ram[23][31:0] = 32'd355283432;
        ram[23][63:32] = 32'd1228061459;
        ram[23][95:64] = 32'd3836173812;
        ram[23][127:96] = 32'd650376785;
        ram[24][31:0] = 32'd1615274362;
        ram[24][63:32] = 32'd3946323928;
        ram[24][95:64] = 32'd2576532341;
        ram[24][127:96] = 32'd3402368761;
        ram[25][31:0] = 32'd3518544175;
        ram[25][63:32] = 32'd2796895359;
        ram[25][95:64] = 32'd457023927;
        ram[25][127:96] = 32'd4006048603;
        ram[26][31:0] = 32'd3745214105;
        ram[26][63:32] = 32'd3574643393;
        ram[26][95:64] = 32'd4071584875;
        ram[26][127:96] = 32'd3862762663;
        ram[27][31:0] = 32'd2414169125;
        ram[27][63:32] = 32'd744992370;
        ram[27][95:64] = 32'd1277603101;
        ram[27][127:96] = 32'd1452439021;
        ram[28][31:0] = 32'd338946051;
        ram[28][63:32] = 32'd958838625;
        ram[28][95:64] = 32'd469884127;
        ram[28][127:96] = 32'd1652892941;
        ram[29][31:0] = 32'd3804836444;
        ram[29][63:32] = 32'd4220214550;
        ram[29][95:64] = 32'd3870599432;
        ram[29][127:96] = 32'd1527611154;
        ram[30][31:0] = 32'd2264552573;
        ram[30][63:32] = 32'd2605200182;
        ram[30][95:64] = 32'd3622924683;
        ram[30][127:96] = 32'd1887842932;
        ram[31][31:0] = 32'd1576649343;
        ram[31][63:32] = 32'd1528221139;
        ram[31][95:64] = 32'd1640972091;
        ram[31][127:96] = 32'd2531376941;
        ram[32][31:0] = 32'd4248669786;
        ram[32][63:32] = 32'd4156816041;
        ram[32][95:64] = 32'd3185392084;
        ram[32][127:96] = 32'd2412978687;
        ram[33][31:0] = 32'd347320602;
        ram[33][63:32] = 32'd1632895041;
        ram[33][95:64] = 32'd3657150815;
        ram[33][127:96] = 32'd1710980134;
        ram[34][31:0] = 32'd3179925528;
        ram[34][63:32] = 32'd3516062355;
        ram[34][95:64] = 32'd1254375529;
        ram[34][127:96] = 32'd1055727677;
        ram[35][31:0] = 32'd452007419;
        ram[35][63:32] = 32'd3732737218;
        ram[35][95:64] = 32'd1891504155;
        ram[35][127:96] = 32'd1991012920;
        ram[36][31:0] = 32'd1650381935;
        ram[36][63:32] = 32'd2063066909;
        ram[36][95:64] = 32'd2237304365;
        ram[36][127:96] = 32'd3636918211;
        ram[37][31:0] = 32'd4188531896;
        ram[37][63:32] = 32'd2114575800;
        ram[37][95:64] = 32'd2984452783;
        ram[37][127:96] = 32'd1108166826;
        ram[38][31:0] = 32'd2253932096;
        ram[38][63:32] = 32'd3061874645;
        ram[38][95:64] = 32'd1372006202;
        ram[38][127:96] = 32'd1567660096;
        ram[39][31:0] = 32'd1564620619;
        ram[39][63:32] = 32'd2310668724;
        ram[39][95:64] = 32'd16933433;
        ram[39][127:96] = 32'd3037698070;
        ram[40][31:0] = 32'd2288570994;
        ram[40][63:32] = 32'd2556436400;
        ram[40][95:64] = 32'd3143417896;
        ram[40][127:96] = 32'd3528470030;
        ram[41][31:0] = 32'd342696692;
        ram[41][63:32] = 32'd3961919093;
        ram[41][95:64] = 32'd2253906058;
        ram[41][127:96] = 32'd367704174;
        ram[42][31:0] = 32'd1042391242;
        ram[42][63:32] = 32'd705866065;
        ram[42][95:64] = 32'd911045719;
        ram[42][127:96] = 32'd4210643370;
        ram[43][31:0] = 32'd3645680872;
        ram[43][63:32] = 32'd1258215212;
        ram[43][95:64] = 32'd2579075201;
        ram[43][127:96] = 32'd3285653861;
        ram[44][31:0] = 32'd563464194;
        ram[44][63:32] = 32'd4089579967;
        ram[44][95:64] = 32'd4072800167;
        ram[44][127:96] = 32'd487094244;
        ram[45][31:0] = 32'd1185846637;
        ram[45][63:32] = 32'd500375006;
        ram[45][95:64] = 32'd3172527317;
        ram[45][127:96] = 32'd1977938445;
        ram[46][31:0] = 32'd424689813;
        ram[46][63:32] = 32'd22147021;
        ram[46][95:64] = 32'd3062031139;
        ram[46][127:96] = 32'd793217816;
        ram[47][31:0] = 32'd2553602888;
        ram[47][63:32] = 32'd669715075;
        ram[47][95:64] = 32'd1502392286;
        ram[47][127:96] = 32'd330133115;
        ram[48][31:0] = 32'd4135019198;
        ram[48][63:32] = 32'd1033777528;
        ram[48][95:64] = 32'd2955644450;
        ram[48][127:96] = 32'd2443887426;
        ram[49][31:0] = 32'd2584950764;
        ram[49][63:32] = 32'd1696743885;
        ram[49][95:64] = 32'd2875093575;
        ram[49][127:96] = 32'd4120401195;
        ram[50][31:0] = 32'd839720366;
        ram[50][63:32] = 32'd3316635280;
        ram[50][95:64] = 32'd538073080;
        ram[50][127:96] = 32'd1831871360;
        ram[51][31:0] = 32'd1535612339;
        ram[51][63:32] = 32'd1390670909;
        ram[51][95:64] = 32'd4213338333;
        ram[51][127:96] = 32'd513445133;
        ram[52][31:0] = 32'd3472524183;
        ram[52][63:32] = 32'd1304622152;
        ram[52][95:64] = 32'd118596569;
        ram[52][127:96] = 32'd4202191155;
        ram[53][31:0] = 32'd2809482033;
        ram[53][63:32] = 32'd4065612688;
        ram[53][95:64] = 32'd635033231;
        ram[53][127:96] = 32'd4098659685;
        ram[54][31:0] = 32'd4112074439;
        ram[54][63:32] = 32'd2718828492;
        ram[54][95:64] = 32'd1056999408;
        ram[54][127:96] = 32'd193565387;
        ram[55][31:0] = 32'd273442298;
        ram[55][63:32] = 32'd3019464660;
        ram[55][95:64] = 32'd1384897455;
        ram[55][127:96] = 32'd408571269;
        ram[56][31:0] = 32'd463140193;
        ram[56][63:32] = 32'd4258929245;
        ram[56][95:64] = 32'd2717548623;
        ram[56][127:96] = 32'd2688484918;
        ram[57][31:0] = 32'd4120475529;
        ram[57][63:32] = 32'd665005425;
        ram[57][95:64] = 32'd2766110621;
        ram[57][127:96] = 32'd2346487764;
        ram[58][31:0] = 32'd3044665406;
        ram[58][63:32] = 32'd2492348860;
        ram[58][95:64] = 32'd3059098805;
        ram[58][127:96] = 32'd379016448;
        ram[59][31:0] = 32'd1954450839;
        ram[59][63:32] = 32'd3293190254;
        ram[59][95:64] = 32'd245166882;
        ram[59][127:96] = 32'd1677771600;
        ram[60][31:0] = 32'd524685732;
        ram[60][63:32] = 32'd3112036660;
        ram[60][95:64] = 32'd502196391;
        ram[60][127:96] = 32'd1440318250;
        ram[61][31:0] = 32'd1318439210;
        ram[61][63:32] = 32'd2541699711;
        ram[61][95:64] = 32'd801919684;
        ram[61][127:96] = 32'd3793934249;
        ram[62][31:0] = 32'd995719055;
        ram[62][63:32] = 32'd3927970277;
        ram[62][95:64] = 32'd3899655140;
        ram[62][127:96] = 32'd3445548488;
        ram[63][31:0] = 32'd2967320824;
        ram[63][63:32] = 32'd2885822038;
        ram[63][95:64] = 32'd2317459088;
        ram[63][127:96] = 32'd3493356248;
        ram[64][31:0] = 32'd2441338571;
        ram[64][63:32] = 32'd3530939413;
        ram[64][95:64] = 32'd1644063503;
        ram[64][127:96] = 32'd1637175110;
        ram[65][31:0] = 32'd1884041322;
        ram[65][63:32] = 32'd1776590124;
        ram[65][95:64] = 32'd2158457297;
        ram[65][127:96] = 32'd2617758261;
        ram[66][31:0] = 32'd4124826968;
        ram[66][63:32] = 32'd2848828629;
        ram[66][95:64] = 32'd2745001205;
        ram[66][127:96] = 32'd2501490696;
        ram[67][31:0] = 32'd2441997828;
        ram[67][63:32] = 32'd90054363;
        ram[67][95:64] = 32'd4155868294;
        ram[67][127:96] = 32'd1009868606;
        ram[68][31:0] = 32'd430353697;
        ram[68][63:32] = 32'd3917527697;
        ram[68][95:64] = 32'd3059870078;
        ram[68][127:96] = 32'd2653768591;
        ram[69][31:0] = 32'd3997787016;
        ram[69][63:32] = 32'd2967447291;
        ram[69][95:64] = 32'd1532905441;
        ram[69][127:96] = 32'd568574415;
        ram[70][31:0] = 32'd469901265;
        ram[70][63:32] = 32'd3708121482;
        ram[70][95:64] = 32'd1881898418;
        ram[70][127:96] = 32'd2307617241;
        ram[71][31:0] = 32'd935136977;
        ram[71][63:32] = 32'd3139190243;
        ram[71][95:64] = 32'd2132904872;
        ram[71][127:96] = 32'd4288613521;
        ram[72][31:0] = 32'd2458363594;
        ram[72][63:32] = 32'd4124324693;
        ram[72][95:64] = 32'd3645826661;
        ram[72][127:96] = 32'd2507289981;
        ram[73][31:0] = 32'd1640016259;
        ram[73][63:32] = 32'd1249044169;
        ram[73][95:64] = 32'd3223530803;
        ram[73][127:96] = 32'd1478684809;
        ram[74][31:0] = 32'd3937584621;
        ram[74][63:32] = 32'd2331663310;
        ram[74][95:64] = 32'd3323657135;
        ram[74][127:96] = 32'd2571156935;
        ram[75][31:0] = 32'd3281353580;
        ram[75][63:32] = 32'd582366332;
        ram[75][95:64] = 32'd3424128274;
        ram[75][127:96] = 32'd4080236004;
        ram[76][31:0] = 32'd800561686;
        ram[76][63:32] = 32'd405757788;
        ram[76][95:64] = 32'd3900608396;
        ram[76][127:96] = 32'd4032726540;
        ram[77][31:0] = 32'd845367245;
        ram[77][63:32] = 32'd1432220972;
        ram[77][95:64] = 32'd727353973;
        ram[77][127:96] = 32'd261335557;
        ram[78][31:0] = 32'd2830282665;
        ram[78][63:32] = 32'd4174569149;
        ram[78][95:64] = 32'd303175971;
        ram[78][127:96] = 32'd735135208;
        ram[79][31:0] = 32'd2596268729;
        ram[79][63:32] = 32'd2714230834;
        ram[79][95:64] = 32'd2835077050;
        ram[79][127:96] = 32'd1482942463;
        ram[80][31:0] = 32'd2364460379;
        ram[80][63:32] = 32'd896564245;
        ram[80][95:64] = 32'd2089037115;
        ram[80][127:96] = 32'd1861217836;
        ram[81][31:0] = 32'd3987095755;
        ram[81][63:32] = 32'd1715720789;
        ram[81][95:64] = 32'd3602797429;
        ram[81][127:96] = 32'd310070123;
        ram[82][31:0] = 32'd77460711;
        ram[82][63:32] = 32'd1741242015;
        ram[82][95:64] = 32'd3508612389;
        ram[82][127:96] = 32'd3184438248;
        ram[83][31:0] = 32'd4266769130;
        ram[83][63:32] = 32'd2296982685;
        ram[83][95:64] = 32'd2783766917;
        ram[83][127:96] = 32'd1195626943;
        ram[84][31:0] = 32'd1688024943;
        ram[84][63:32] = 32'd3322552394;
        ram[84][95:64] = 32'd1821314294;
        ram[84][127:96] = 32'd3023854751;
        ram[85][31:0] = 32'd1638179589;
        ram[85][63:32] = 32'd315843574;
        ram[85][95:64] = 32'd3024089183;
        ram[85][127:96] = 32'd2846218665;
        ram[86][31:0] = 32'd1668394988;
        ram[86][63:32] = 32'd2791959723;
        ram[86][95:64] = 32'd3770003965;
        ram[86][127:96] = 32'd4150740891;
        ram[87][31:0] = 32'd904943400;
        ram[87][63:32] = 32'd3103175904;
        ram[87][95:64] = 32'd1182201995;
        ram[87][127:96] = 32'd2365388450;
        ram[88][31:0] = 32'd163922335;
        ram[88][63:32] = 32'd3565100911;
        ram[88][95:64] = 32'd2972176425;
        ram[88][127:96] = 32'd3917761171;
        ram[89][31:0] = 32'd2257235136;
        ram[89][63:32] = 32'd3927443995;
        ram[89][95:64] = 32'd3685422029;
        ram[89][127:96] = 32'd3154057553;
        ram[90][31:0] = 32'd3069921140;
        ram[90][63:32] = 32'd3378581894;
        ram[90][95:64] = 32'd2935077560;
        ram[90][127:96] = 32'd2723076636;
        ram[91][31:0] = 32'd1333182938;
        ram[91][63:32] = 32'd1161783265;
        ram[91][95:64] = 32'd2025896452;
        ram[91][127:96] = 32'd1351470440;
        ram[92][31:0] = 32'd4078620521;
        ram[92][63:32] = 32'd2305103248;
        ram[92][95:64] = 32'd4146930610;
        ram[92][127:96] = 32'd2775974076;
        ram[93][31:0] = 32'd3653485486;
        ram[93][63:32] = 32'd3628187523;
        ram[93][95:64] = 32'd2971708932;
        ram[93][127:96] = 32'd2719622023;
        ram[94][31:0] = 32'd3828805185;
        ram[94][63:32] = 32'd436835430;
        ram[94][95:64] = 32'd515798227;
        ram[94][127:96] = 32'd708784957;
        ram[95][31:0] = 32'd1150466899;
        ram[95][63:32] = 32'd1741094807;
        ram[95][95:64] = 32'd3223401649;
        ram[95][127:96] = 32'd636051292;
        ram[96][31:0] = 32'd3274611019;
        ram[96][63:32] = 32'd817202464;
        ram[96][95:64] = 32'd1481982667;
        ram[96][127:96] = 32'd4132411223;
        ram[97][31:0] = 32'd3781905541;
        ram[97][63:32] = 32'd3497432784;
        ram[97][95:64] = 32'd2210144971;
        ram[97][127:96] = 32'd3183432554;
        ram[98][31:0] = 32'd2117412331;
        ram[98][63:32] = 32'd479449245;
        ram[98][95:64] = 32'd1469178574;
        ram[98][127:96] = 32'd1515244782;
        ram[99][31:0] = 32'd3733634737;
        ram[99][63:32] = 32'd353205820;
        ram[99][95:64] = 32'd3505084960;
        ram[99][127:96] = 32'd509805444;
        ram[100][31:0] = 32'd2244076081;
        ram[100][63:32] = 32'd427139017;
        ram[100][95:64] = 32'd2447482056;
        ram[100][127:96] = 32'd3705260287;
        ram[101][31:0] = 32'd602052412;
        ram[101][63:32] = 32'd1195841942;
        ram[101][95:64] = 32'd532774694;
        ram[101][127:96] = 32'd4228653296;
        ram[102][31:0] = 32'd1991242564;
        ram[102][63:32] = 32'd881702054;
        ram[102][95:64] = 32'd3442998655;
        ram[102][127:96] = 32'd2509072348;
        ram[103][31:0] = 32'd3063633923;
        ram[103][63:32] = 32'd4263007220;
        ram[103][95:64] = 32'd2622463751;
        ram[103][127:96] = 32'd2483981373;
        ram[104][31:0] = 32'd3762483973;
        ram[104][63:32] = 32'd857483597;
        ram[104][95:64] = 32'd3304050455;
        ram[104][127:96] = 32'd3868382538;
        ram[105][31:0] = 32'd2008269494;
        ram[105][63:32] = 32'd3124744987;
        ram[105][95:64] = 32'd2139306794;
        ram[105][127:96] = 32'd3226229557;
        ram[106][31:0] = 32'd4107482093;
        ram[106][63:32] = 32'd3487355990;
        ram[106][95:64] = 32'd887963095;
        ram[106][127:96] = 32'd1334217002;
        ram[107][31:0] = 32'd807619004;
        ram[107][63:32] = 32'd3047596899;
        ram[107][95:64] = 32'd896214945;
        ram[107][127:96] = 32'd3279784998;
        ram[108][31:0] = 32'd842198295;
        ram[108][63:32] = 32'd816551425;
        ram[108][95:64] = 32'd1408779004;
        ram[108][127:96] = 32'd2315575124;
        ram[109][31:0] = 32'd4034103201;
        ram[109][63:32] = 32'd465935354;
        ram[109][95:64] = 32'd636048466;
        ram[109][127:96] = 32'd2807691332;
        ram[110][31:0] = 32'd3456116014;
        ram[110][63:32] = 32'd924466934;
        ram[110][95:64] = 32'd2950643337;
        ram[110][127:96] = 32'd1586603011;
        ram[111][31:0] = 32'd2677223067;
        ram[111][63:32] = 32'd3509235017;
        ram[111][95:64] = 32'd1320511667;
        ram[111][127:96] = 32'd3084548448;
        ram[112][31:0] = 32'd2047532963;
        ram[112][63:32] = 32'd658651725;
        ram[112][95:64] = 32'd2853006304;
        ram[112][127:96] = 32'd201021719;
        ram[113][31:0] = 32'd1012981055;
        ram[113][63:32] = 32'd4144249236;
        ram[113][95:64] = 32'd1488664850;
        ram[113][127:96] = 32'd4791580;
        ram[114][31:0] = 32'd2010861474;
        ram[114][63:32] = 32'd96864288;
        ram[114][95:64] = 32'd4143306261;
        ram[114][127:96] = 32'd1894780540;
        ram[115][31:0] = 32'd334824474;
        ram[115][63:32] = 32'd2515252354;
        ram[115][95:64] = 32'd2318869365;
        ram[115][127:96] = 32'd909928079;
        ram[116][31:0] = 32'd3521762258;
        ram[116][63:32] = 32'd1435079633;
        ram[116][95:64] = 32'd2321964682;
        ram[116][127:96] = 32'd1444845120;
        ram[117][31:0] = 32'd3544189000;
        ram[117][63:32] = 32'd821820080;
        ram[117][95:64] = 32'd1889226206;
        ram[117][127:96] = 32'd2169217366;
        ram[118][31:0] = 32'd1119598195;
        ram[118][63:32] = 32'd4114965494;
        ram[118][95:64] = 32'd2841812471;
        ram[118][127:96] = 32'd3061835182;
        ram[119][31:0] = 32'd1839489904;
        ram[119][63:32] = 32'd815049655;
        ram[119][95:64] = 32'd2289392119;
        ram[119][127:96] = 32'd840506018;
        ram[120][31:0] = 32'd125390000;
        ram[120][63:32] = 32'd2639408353;
        ram[120][95:64] = 32'd3393357937;
        ram[120][127:96] = 32'd3327007420;
        ram[121][31:0] = 32'd998179708;
        ram[121][63:32] = 32'd1497784997;
        ram[121][95:64] = 32'd3551446877;
        ram[121][127:96] = 32'd1179387712;
        ram[122][31:0] = 32'd3230286556;
        ram[122][63:32] = 32'd654573334;
        ram[122][95:64] = 32'd4090258182;
        ram[122][127:96] = 32'd2199790567;
        ram[123][31:0] = 32'd2583156540;
        ram[123][63:32] = 32'd2115438628;
        ram[123][95:64] = 32'd4244092772;
        ram[123][127:96] = 32'd1834135079;
        ram[124][31:0] = 32'd863026729;
        ram[124][63:32] = 32'd3663618438;
        ram[124][95:64] = 32'd4163492510;
        ram[124][127:96] = 32'd1344952170;
        ram[125][31:0] = 32'd3426938455;
        ram[125][63:32] = 32'd2592532499;
        ram[125][95:64] = 32'd1661402023;
        ram[125][127:96] = 32'd1431025879;
        ram[126][31:0] = 32'd225331988;
        ram[126][63:32] = 32'd3200330407;
        ram[126][95:64] = 32'd4068327518;
        ram[126][127:96] = 32'd3984605869;
        ram[127][31:0] = 32'd1247575968;
        ram[127][63:32] = 32'd1995849586;
        ram[127][95:64] = 32'd513403764;
        ram[127][127:96] = 32'd4030006546;
        ram[128][31:0] = 32'd1581423827;
        ram[128][63:32] = 32'd421452164;
        ram[128][95:64] = 32'd2973446334;
        ram[128][127:96] = 32'd4209937496;
        ram[129][31:0] = 32'd1918061132;
        ram[129][63:32] = 32'd4067077614;
        ram[129][95:64] = 32'd849664853;
        ram[129][127:96] = 32'd1902800231;
        ram[130][31:0] = 32'd2563473161;
        ram[130][63:32] = 32'd3220870596;
        ram[130][95:64] = 32'd3048636483;
        ram[130][127:96] = 32'd2950126546;
        ram[131][31:0] = 32'd1326168490;
        ram[131][63:32] = 32'd1316917817;
        ram[131][95:64] = 32'd736640889;
        ram[131][127:96] = 32'd3884199812;
        ram[132][31:0] = 32'd4183271945;
        ram[132][63:32] = 32'd730554504;
        ram[132][95:64] = 32'd1157531596;
        ram[132][127:96] = 32'd3014035020;
        ram[133][31:0] = 32'd1996478713;
        ram[133][63:32] = 32'd1603575421;
        ram[133][95:64] = 32'd2544290285;
        ram[133][127:96] = 32'd1551618470;
        ram[134][31:0] = 32'd4216548472;
        ram[134][63:32] = 32'd1269482248;
        ram[134][95:64] = 32'd2662158238;
        ram[134][127:96] = 32'd1252831804;
        ram[135][31:0] = 32'd3769408227;
        ram[135][63:32] = 32'd3630666215;
        ram[135][95:64] = 32'd2523859335;
        ram[135][127:96] = 32'd108826463;
        ram[136][31:0] = 32'd3265468743;
        ram[136][63:32] = 32'd3521037345;
        ram[136][95:64] = 32'd3953366411;
        ram[136][127:96] = 32'd1615745349;
        ram[137][31:0] = 32'd924290257;
        ram[137][63:32] = 32'd3932271196;
        ram[137][95:64] = 32'd828402464;
        ram[137][127:96] = 32'd3755615061;
        ram[138][31:0] = 32'd2229852656;
        ram[138][63:32] = 32'd3462769718;
        ram[138][95:64] = 32'd1152867193;
        ram[138][127:96] = 32'd3459416445;
        ram[139][31:0] = 32'd2229379164;
        ram[139][63:32] = 32'd2146319491;
        ram[139][95:64] = 32'd1593008829;
        ram[139][127:96] = 32'd1691044550;
        ram[140][31:0] = 32'd2338900121;
        ram[140][63:32] = 32'd2094957369;
        ram[140][95:64] = 32'd3011983409;
        ram[140][127:96] = 32'd3434699751;
        ram[141][31:0] = 32'd869541130;
        ram[141][63:32] = 32'd1601476386;
        ram[141][95:64] = 32'd1705309202;
        ram[141][127:96] = 32'd1925411768;
        ram[142][31:0] = 32'd1475611248;
        ram[142][63:32] = 32'd3732094373;
        ram[142][95:64] = 32'd4180903970;
        ram[142][127:96] = 32'd533451981;
        ram[143][31:0] = 32'd403146832;
        ram[143][63:32] = 32'd660266423;
        ram[143][95:64] = 32'd4096603703;
        ram[143][127:96] = 32'd522515645;
        ram[144][31:0] = 32'd1716076338;
        ram[144][63:32] = 32'd469589016;
        ram[144][95:64] = 32'd3176129940;
        ram[144][127:96] = 32'd2815817156;
        ram[145][31:0] = 32'd914006725;
        ram[145][63:32] = 32'd483805297;
        ram[145][95:64] = 32'd1239020060;
        ram[145][127:96] = 32'd3440524923;
        ram[146][31:0] = 32'd3939647983;
        ram[146][63:32] = 32'd1423656890;
        ram[146][95:64] = 32'd2066734253;
        ram[146][127:96] = 32'd1101126375;
        ram[147][31:0] = 32'd3233337789;
        ram[147][63:32] = 32'd2182645025;
        ram[147][95:64] = 32'd403378138;
        ram[147][127:96] = 32'd1386873771;
        ram[148][31:0] = 32'd2408379302;
        ram[148][63:32] = 32'd2126572521;
        ram[148][95:64] = 32'd3082553007;
        ram[148][127:96] = 32'd1646515767;
        ram[149][31:0] = 32'd2888243094;
        ram[149][63:32] = 32'd3535940700;
        ram[149][95:64] = 32'd218926266;
        ram[149][127:96] = 32'd699313956;
        ram[150][31:0] = 32'd699365697;
        ram[150][63:32] = 32'd1061024359;
        ram[150][95:64] = 32'd523974119;
        ram[150][127:96] = 32'd1949152991;
        ram[151][31:0] = 32'd4057563322;
        ram[151][63:32] = 32'd1618144234;
        ram[151][95:64] = 32'd920782161;
        ram[151][127:96] = 32'd3986635328;
        ram[152][31:0] = 32'd2953791377;
        ram[152][63:32] = 32'd3511563354;
        ram[152][95:64] = 32'd2559326217;
        ram[152][127:96] = 32'd160596143;
        ram[153][31:0] = 32'd702302819;
        ram[153][63:32] = 32'd600314913;
        ram[153][95:64] = 32'd1036899548;
        ram[153][127:96] = 32'd4288664088;
        ram[154][31:0] = 32'd3292421464;
        ram[154][63:32] = 32'd1266899086;
        ram[154][95:64] = 32'd3524599878;
        ram[154][127:96] = 32'd11211046;
        ram[155][31:0] = 32'd2147528937;
        ram[155][63:32] = 32'd765391404;
        ram[155][95:64] = 32'd650152461;
        ram[155][127:96] = 32'd2373385250;
        ram[156][31:0] = 32'd3691275069;
        ram[156][63:32] = 32'd1909344899;
        ram[156][95:64] = 32'd3411209394;
        ram[156][127:96] = 32'd111369000;
        ram[157][31:0] = 32'd108823116;
        ram[157][63:32] = 32'd4225840529;
        ram[157][95:64] = 32'd911457724;
        ram[157][127:96] = 32'd4116914749;
        ram[158][31:0] = 32'd86211075;
        ram[158][63:32] = 32'd1090431518;
        ram[158][95:64] = 32'd3651902078;
        ram[158][127:96] = 32'd3605989952;
        ram[159][31:0] = 32'd1543105877;
        ram[159][63:32] = 32'd107830373;
        ram[159][95:64] = 32'd3568991821;
        ram[159][127:96] = 32'd3147882387;
        ram[160][31:0] = 32'd3889086438;
        ram[160][63:32] = 32'd3812820741;
        ram[160][95:64] = 32'd1424094667;
        ram[160][127:96] = 32'd4067317687;
        ram[161][31:0] = 32'd550544246;
        ram[161][63:32] = 32'd1749328043;
        ram[161][95:64] = 32'd1276954913;
        ram[161][127:96] = 32'd2034393425;
        ram[162][31:0] = 32'd2300180881;
        ram[162][63:32] = 32'd4206062990;
        ram[162][95:64] = 32'd2784853932;
        ram[162][127:96] = 32'd322357615;
        ram[163][31:0] = 32'd2701092793;
        ram[163][63:32] = 32'd1452550502;
        ram[163][95:64] = 32'd3786347631;
        ram[163][127:96] = 32'd2522894847;
        ram[164][31:0] = 32'd2873453145;
        ram[164][63:32] = 32'd2813359384;
        ram[164][95:64] = 32'd3120144388;
        ram[164][127:96] = 32'd475659489;
        ram[165][31:0] = 32'd1936867947;
        ram[165][63:32] = 32'd3080712060;
        ram[165][95:64] = 32'd4159685436;
        ram[165][127:96] = 32'd89312420;
        ram[166][31:0] = 32'd4123313617;
        ram[166][63:32] = 32'd3823881563;
        ram[166][95:64] = 32'd812647693;
        ram[166][127:96] = 32'd560999711;
        ram[167][31:0] = 32'd4073128129;
        ram[167][63:32] = 32'd716422625;
        ram[167][95:64] = 32'd606154580;
        ram[167][127:96] = 32'd2151985146;
        ram[168][31:0] = 32'd2072267703;
        ram[168][63:32] = 32'd2206060871;
        ram[168][95:64] = 32'd1911503576;
        ram[168][127:96] = 32'd3430516374;
        ram[169][31:0] = 32'd662578081;
        ram[169][63:32] = 32'd2331235146;
        ram[169][95:64] = 32'd899706535;
        ram[169][127:96] = 32'd528435148;
        ram[170][31:0] = 32'd772379733;
        ram[170][63:32] = 32'd85007220;
        ram[170][95:64] = 32'd666405120;
        ram[170][127:96] = 32'd1731237928;
        ram[171][31:0] = 32'd781313041;
        ram[171][63:32] = 32'd1329909483;
        ram[171][95:64] = 32'd4109187007;
        ram[171][127:96] = 32'd1220117427;
        ram[172][31:0] = 32'd2293783707;
        ram[172][63:32] = 32'd2765668052;
        ram[172][95:64] = 32'd1050749044;
        ram[172][127:96] = 32'd168821635;
        ram[173][31:0] = 32'd984956215;
        ram[173][63:32] = 32'd1341386525;
        ram[173][95:64] = 32'd3300358697;
        ram[173][127:96] = 32'd4204941700;
        ram[174][31:0] = 32'd2824012066;
        ram[174][63:32] = 32'd2908751719;
        ram[174][95:64] = 32'd2093503010;
        ram[174][127:96] = 32'd3070843493;
        ram[175][31:0] = 32'd1020382117;
        ram[175][63:32] = 32'd440612704;
        ram[175][95:64] = 32'd1945165593;
        ram[175][127:96] = 32'd2023405860;
        ram[176][31:0] = 32'd266762623;
        ram[176][63:32] = 32'd76247026;
        ram[176][95:64] = 32'd3602815316;
        ram[176][127:96] = 32'd3409958362;
        ram[177][31:0] = 32'd3004227477;
        ram[177][63:32] = 32'd265858089;
        ram[177][95:64] = 32'd2490057219;
        ram[177][127:96] = 32'd2444809984;
        ram[178][31:0] = 32'd265621438;
        ram[178][63:32] = 32'd3501601674;
        ram[178][95:64] = 32'd299549045;
        ram[178][127:96] = 32'd3297497505;
        ram[179][31:0] = 32'd292650974;
        ram[179][63:32] = 32'd2752499399;
        ram[179][95:64] = 32'd3656605274;
        ram[179][127:96] = 32'd602760059;
        ram[180][31:0] = 32'd264781874;
        ram[180][63:32] = 32'd3453091153;
        ram[180][95:64] = 32'd1583494039;
        ram[180][127:96] = 32'd2532020940;
        ram[181][31:0] = 32'd1061855659;
        ram[181][63:32] = 32'd137891339;
        ram[181][95:64] = 32'd2075556532;
        ram[181][127:96] = 32'd2678040300;
        ram[182][31:0] = 32'd69884107;
        ram[182][63:32] = 32'd1439363931;
        ram[182][95:64] = 32'd2998442618;
        ram[182][127:96] = 32'd3605685312;
        ram[183][31:0] = 32'd1766000469;
        ram[183][63:32] = 32'd3548136803;
        ram[183][95:64] = 32'd3288289380;
        ram[183][127:96] = 32'd27263033;
        ram[184][31:0] = 32'd3833161201;
        ram[184][63:32] = 32'd2458406238;
        ram[184][95:64] = 32'd162191551;
        ram[184][127:96] = 32'd2692232349;
        ram[185][31:0] = 32'd725439312;
        ram[185][63:32] = 32'd336889000;
        ram[185][95:64] = 32'd3311420871;
        ram[185][127:96] = 32'd3044130341;
        ram[186][31:0] = 32'd1292464610;
        ram[186][63:32] = 32'd4084688614;
        ram[186][95:64] = 32'd689947192;
        ram[186][127:96] = 32'd2111772806;
        ram[187][31:0] = 32'd292433743;
        ram[187][63:32] = 32'd821619415;
        ram[187][95:64] = 32'd1056728340;
        ram[187][127:96] = 32'd811162109;
        ram[188][31:0] = 32'd3332007732;
        ram[188][63:32] = 32'd857701527;
        ram[188][95:64] = 32'd1731907904;
        ram[188][127:96] = 32'd1320792984;
        ram[189][31:0] = 32'd2829182134;
        ram[189][63:32] = 32'd2869663792;
        ram[189][95:64] = 32'd3678702924;
        ram[189][127:96] = 32'd3506733921;
        ram[190][31:0] = 32'd3222496793;
        ram[190][63:32] = 32'd813817359;
        ram[190][95:64] = 32'd991043089;
        ram[190][127:96] = 32'd407903955;
        ram[191][31:0] = 32'd909334423;
        ram[191][63:32] = 32'd3599204608;
        ram[191][95:64] = 32'd163370680;
        ram[191][127:96] = 32'd51594790;
        ram[192][31:0] = 32'd2995316459;
        ram[192][63:32] = 32'd2466504171;
        ram[192][95:64] = 32'd1650901911;
        ram[192][127:96] = 32'd3324619571;
        ram[193][31:0] = 32'd1354814296;
        ram[193][63:32] = 32'd2757463226;
        ram[193][95:64] = 32'd3061105897;
        ram[193][127:96] = 32'd2078638802;
        ram[194][31:0] = 32'd3351180924;
        ram[194][63:32] = 32'd2415931644;
        ram[194][95:64] = 32'd840840300;
        ram[194][127:96] = 32'd1735230795;
        ram[195][31:0] = 32'd1340653029;
        ram[195][63:32] = 32'd3010039094;
        ram[195][95:64] = 32'd4291708288;
        ram[195][127:96] = 32'd655375125;
        ram[196][31:0] = 32'd2528156350;
        ram[196][63:32] = 32'd2189076806;
        ram[196][95:64] = 32'd4292686456;
        ram[196][127:96] = 32'd1435160092;
        ram[197][31:0] = 32'd3967436273;
        ram[197][63:32] = 32'd1888095334;
        ram[197][95:64] = 32'd2157703382;
        ram[197][127:96] = 32'd1151411794;
        ram[198][31:0] = 32'd2314760705;
        ram[198][63:32] = 32'd760744189;
        ram[198][95:64] = 32'd329858931;
        ram[198][127:96] = 32'd2128607902;
        ram[199][31:0] = 32'd4275211649;
        ram[199][63:32] = 32'd115316762;
        ram[199][95:64] = 32'd4098353399;
        ram[199][127:96] = 32'd2572948599;
        ram[200][31:0] = 32'd754500382;
        ram[200][63:32] = 32'd3939763522;
        ram[200][95:64] = 32'd3959741461;
        ram[200][127:96] = 32'd2717076327;
        ram[201][31:0] = 32'd3891346024;
        ram[201][63:32] = 32'd571201105;
        ram[201][95:64] = 32'd3027734468;
        ram[201][127:96] = 32'd765267270;
        ram[202][31:0] = 32'd158874295;
        ram[202][63:32] = 32'd756026935;
        ram[202][95:64] = 32'd4071171221;
        ram[202][127:96] = 32'd2606956921;
        ram[203][31:0] = 32'd1965390572;
        ram[203][63:32] = 32'd3131080877;
        ram[203][95:64] = 32'd2532614522;
        ram[203][127:96] = 32'd116081840;
        ram[204][31:0] = 32'd2089907260;
        ram[204][63:32] = 32'd4290118485;
        ram[204][95:64] = 32'd1746275809;
        ram[204][127:96] = 32'd196757670;
        ram[205][31:0] = 32'd3200758228;
        ram[205][63:32] = 32'd959016053;
        ram[205][95:64] = 32'd2790105153;
        ram[205][127:96] = 32'd2118102746;
        ram[206][31:0] = 32'd4185437212;
        ram[206][63:32] = 32'd1444494147;
        ram[206][95:64] = 32'd1698091505;
        ram[206][127:96] = 32'd4271161680;
        ram[207][31:0] = 32'd3143336390;
        ram[207][63:32] = 32'd2471067861;
        ram[207][95:64] = 32'd2151514164;
        ram[207][127:96] = 32'd3512387836;
        ram[208][31:0] = 32'd2442866266;
        ram[208][63:32] = 32'd807590553;
        ram[208][95:64] = 32'd1624961981;
        ram[208][127:96] = 32'd3185900460;
        ram[209][31:0] = 32'd2868439311;
        ram[209][63:32] = 32'd2522320532;
        ram[209][95:64] = 32'd2598268969;
        ram[209][127:96] = 32'd2544945082;
        ram[210][31:0] = 32'd2690967453;
        ram[210][63:32] = 32'd3495259579;
        ram[210][95:64] = 32'd1301565224;
        ram[210][127:96] = 32'd3444648562;
        ram[211][31:0] = 32'd1540859185;
        ram[211][63:32] = 32'd2710526860;
        ram[211][95:64] = 32'd3129315442;
        ram[211][127:96] = 32'd1929108195;
        ram[212][31:0] = 32'd2055262394;
        ram[212][63:32] = 32'd544467061;
        ram[212][95:64] = 32'd1598966603;
        ram[212][127:96] = 32'd528403755;
        ram[213][31:0] = 32'd1681580087;
        ram[213][63:32] = 32'd1560350512;
        ram[213][95:64] = 32'd2265029546;
        ram[213][127:96] = 32'd325563839;
        ram[214][31:0] = 32'd1518218722;
        ram[214][63:32] = 32'd456204038;
        ram[214][95:64] = 32'd2316112060;
        ram[214][127:96] = 32'd19128930;
        ram[215][31:0] = 32'd9740189;
        ram[215][63:32] = 32'd3718178245;
        ram[215][95:64] = 32'd1164318928;
        ram[215][127:96] = 32'd3181973309;
        ram[216][31:0] = 32'd2757871746;
        ram[216][63:32] = 32'd2442557656;
        ram[216][95:64] = 32'd864189442;
        ram[216][127:96] = 32'd4191967086;
        ram[217][31:0] = 32'd1517292233;
        ram[217][63:32] = 32'd1232072696;
        ram[217][95:64] = 32'd747559002;
        ram[217][127:96] = 32'd2792938922;
        ram[218][31:0] = 32'd3833194746;
        ram[218][63:32] = 32'd1352952223;
        ram[218][95:64] = 32'd3917285502;
        ram[218][127:96] = 32'd192059718;
        ram[219][31:0] = 32'd3736677355;
        ram[219][63:32] = 32'd596443674;
        ram[219][95:64] = 32'd3420207582;
        ram[219][127:96] = 32'd4085858993;
        ram[220][31:0] = 32'd1009940429;
        ram[220][63:32] = 32'd3579846374;
        ram[220][95:64] = 32'd386405139;
        ram[220][127:96] = 32'd1933304197;
        ram[221][31:0] = 32'd1024624892;
        ram[221][63:32] = 32'd3827515349;
        ram[221][95:64] = 32'd4090995992;
        ram[221][127:96] = 32'd2573163800;
        ram[222][31:0] = 32'd1306365210;
        ram[222][63:32] = 32'd2522291656;
        ram[222][95:64] = 32'd1364501689;
        ram[222][127:96] = 32'd3155621446;
        ram[223][31:0] = 32'd669111840;
        ram[223][63:32] = 32'd278268436;
        ram[223][95:64] = 32'd391382463;
        ram[223][127:96] = 32'd1907386417;
        ram[224][31:0] = 32'd1245387932;
        ram[224][63:32] = 32'd1758044350;
        ram[224][95:64] = 32'd3864664240;
        ram[224][127:96] = 32'd1022507848;
        ram[225][31:0] = 32'd3469687493;
        ram[225][63:32] = 32'd836715634;
        ram[225][95:64] = 32'd517865842;
        ram[225][127:96] = 32'd4202993744;
        ram[226][31:0] = 32'd3478950353;
        ram[226][63:32] = 32'd2018867184;
        ram[226][95:64] = 32'd3998543292;
        ram[226][127:96] = 32'd2173475915;
        ram[227][31:0] = 32'd565450044;
        ram[227][63:32] = 32'd3133805742;
        ram[227][95:64] = 32'd1596033064;
        ram[227][127:96] = 32'd2521923331;
        ram[228][31:0] = 32'd3267133870;
        ram[228][63:32] = 32'd2193415700;
        ram[228][95:64] = 32'd2456895004;
        ram[228][127:96] = 32'd2683310477;
        ram[229][31:0] = 32'd1120736423;
        ram[229][63:32] = 32'd2827507563;
        ram[229][95:64] = 32'd942389263;
        ram[229][127:96] = 32'd3709315097;
        ram[230][31:0] = 32'd2557444003;
        ram[230][63:32] = 32'd3242730381;
        ram[230][95:64] = 32'd1197034866;
        ram[230][127:96] = 32'd2212276299;
        ram[231][31:0] = 32'd3076543218;
        ram[231][63:32] = 32'd3444626246;
        ram[231][95:64] = 32'd726676612;
        ram[231][127:96] = 32'd416978341;
        ram[232][31:0] = 32'd3748561664;
        ram[232][63:32] = 32'd3169898984;
        ram[232][95:64] = 32'd1164254761;
        ram[232][127:96] = 32'd4204922469;
        ram[233][31:0] = 32'd2044109763;
        ram[233][63:32] = 32'd3586314489;
        ram[233][95:64] = 32'd1840334227;
        ram[233][127:96] = 32'd2918620527;
        ram[234][31:0] = 32'd76708806;
        ram[234][63:32] = 32'd1191377286;
        ram[234][95:64] = 32'd3392235772;
        ram[234][127:96] = 32'd775116840;
        ram[235][31:0] = 32'd63193559;
        ram[235][63:32] = 32'd1199592277;
        ram[235][95:64] = 32'd1105141139;
        ram[235][127:96] = 32'd2153687124;
        ram[236][31:0] = 32'd4223266270;
        ram[236][63:32] = 32'd2788157755;
        ram[236][95:64] = 32'd2141896945;
        ram[236][127:96] = 32'd2534706481;
        ram[237][31:0] = 32'd1116008264;
        ram[237][63:32] = 32'd2913893151;
        ram[237][95:64] = 32'd2097728883;
        ram[237][127:96] = 32'd3700264061;
        ram[238][31:0] = 32'd1618745728;
        ram[238][63:32] = 32'd1906659600;
        ram[238][95:64] = 32'd3692314337;
        ram[238][127:96] = 32'd1233392266;
        ram[239][31:0] = 32'd2529817444;
        ram[239][63:32] = 32'd2432425057;
        ram[239][95:64] = 32'd1887635491;
        ram[239][127:96] = 32'd1670570220;
        ram[240][31:0] = 32'd269126776;
        ram[240][63:32] = 32'd1162456992;
        ram[240][95:64] = 32'd706727247;
        ram[240][127:96] = 32'd3714607084;
        ram[241][31:0] = 32'd2358691;
        ram[241][63:32] = 32'd3011036640;
        ram[241][95:64] = 32'd2186720106;
        ram[241][127:96] = 32'd227677533;
        ram[242][31:0] = 32'd1940244178;
        ram[242][63:32] = 32'd1355465943;
        ram[242][95:64] = 32'd2846411311;
        ram[242][127:96] = 32'd1340868090;
        ram[243][31:0] = 32'd3134925533;
        ram[243][63:32] = 32'd2724948106;
        ram[243][95:64] = 32'd3423332702;
        ram[243][127:96] = 32'd267738865;
        ram[244][31:0] = 32'd1273610730;
        ram[244][63:32] = 32'd380731391;
        ram[244][95:64] = 32'd2323391226;
        ram[244][127:96] = 32'd431221963;
        ram[245][31:0] = 32'd3930060900;
        ram[245][63:32] = 32'd2623441966;
        ram[245][95:64] = 32'd2934343038;
        ram[245][127:96] = 32'd1323475681;
        ram[246][31:0] = 32'd2138509856;
        ram[246][63:32] = 32'd957211627;
        ram[246][95:64] = 32'd3822672388;
        ram[246][127:96] = 32'd1952340139;
        ram[247][31:0] = 32'd3995363066;
        ram[247][63:32] = 32'd4181739735;
        ram[247][95:64] = 32'd3997510275;
        ram[247][127:96] = 32'd88478458;
        ram[248][31:0] = 32'd669592020;
        ram[248][63:32] = 32'd1916779651;
        ram[248][95:64] = 32'd532973784;
        ram[248][127:96] = 32'd55503118;
        ram[249][31:0] = 32'd1855610634;
        ram[249][63:32] = 32'd2243105101;
        ram[249][95:64] = 32'd2364278147;
        ram[249][127:96] = 32'd1429796383;
        ram[250][31:0] = 32'd136122382;
        ram[250][63:32] = 32'd1757685921;
        ram[250][95:64] = 32'd1476013580;
        ram[250][127:96] = 32'd1864759393;
        ram[251][31:0] = 32'd2136110024;
        ram[251][63:32] = 32'd2395804748;
        ram[251][95:64] = 32'd479112565;
        ram[251][127:96] = 32'd4059948122;
        ram[252][31:0] = 32'd4049834946;
        ram[252][63:32] = 32'd2905712961;
        ram[252][95:64] = 32'd1079389392;
        ram[252][127:96] = 32'd743506454;
        ram[253][31:0] = 32'd891830012;
        ram[253][63:32] = 32'd354624723;
        ram[253][95:64] = 32'd1182686270;
        ram[253][127:96] = 32'd2560991281;
        ram[254][31:0] = 32'd3935014123;
        ram[254][63:32] = 32'd1703702969;
        ram[254][95:64] = 32'd1682531465;
        ram[254][127:96] = 32'd361342986;
        ram[255][31:0] = 32'd1804380535;
        ram[255][63:32] = 32'd1888120797;
        ram[255][95:64] = 32'd1248002737;
        ram[255][127:96] = 32'd3621827067;

    end
    always @(posedge clk) begin
        addr_r <= raddr;
        if(we) ram[waddr] <= din;
    end
    assign dout = ram[addr_r]; 

endmodule
