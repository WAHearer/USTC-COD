
/*
本文件是一个测试文件，用于测试cache模块
工作原理是模仿CPU的读写请求，对cache进行读写操作
将Cache返回的数据与预先数据进行比较，如果一致则测试通过
*/
`timescale 1ns/1ps
module cache_tb();

    //测试参数
    parameter READ_NUM = 2000;  // 测试次数 这里设置为2000次读，1000次写
    parameter WRITE_NUM = 1000;  
    //模块参数
    parameter INDEX_WIDTH       = 3;   // Cache索引位宽 2^3=8行
    parameter LINE_OFFSET_WIDTH = 2;   // 行偏移位宽，决定了一行的宽度 2^2=4字
    parameter SPACE_OFFSET      = 2;   // 一个地址空间占1个字节，因此一个字需要4个地址空间，由于假设为整字读取，处理地址的时候可以默认后两位为0
    parameter MEM_ADDR_WIDTH    = 10;   // 为了简化，这里假设内存地址宽度为10位（CPU请求地址仍然是32位，只不过我们这里简化处理，截断了高位） 
    parameter WAY_NUM           = 1;   // Cache N路组相联(N=1的时候是直接映射)

    // 变化的信号 CPU发出
    reg clk=1;
    reg rstn=1;
    reg stat=0;
    // 等rstn信号稳定后 clk信号才开始翻转
    initial begin
        #1 rstn = 0;
        #1 rstn = 1;
        stat = 1;
    end
    always  #1 clk = ~clk;

    wire [31:0] addr;
    wire r_req;
    wire w_req;
    wire [31:0] w_data;

    // 导线
    wire [31:0] r_data;
    wire miss;
    wire mem_r;
    wire mem_w;
    wire [31:0] mem_addr;
    wire [127:0] mem_w_data;
    wire [127:0] mem_r_data;
    wire mem_ready;

    // 用于测试的信号
    reg [MEM_ADDR_WIDTH-1:0] test_addr[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试地址
    reg [32:0] test_data[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试数据 最高位用于标记是否写入 0：读 1：写
    reg [31:0] test_cnt=0;  // 用于计数，每次读写操作后加1
    reg diff=0;  // 用于标记是否有不一致的数据

    // 用于对比的提交，当前cache应该给出的数据
    wire op;
    wire[31:0] data;
    assign op = test_data[test_cnt-1][32];
    assign data = test_data[test_cnt-1][31:0];
    
    // 状态机
    assign addr = test_addr[test_cnt]<<SPACE_OFFSET;
    assign r_req = test_data[test_cnt][32] == 0 ? 1 : 0;
    assign w_req = test_data[test_cnt][32] == 1 ? 1 : 0;
    assign w_data = test_data[test_cnt][31:0];
    always @(posedge clk) begin
        if (!miss && (test_cnt < READ_NUM+WRITE_NUM) && stat) begin
            if (test_data[test_cnt-1][32] == 0) begin  // 读
                if (r_data != test_data[test_cnt-1][31:0]) begin
                    $display("Read error at %d, expect %h, get %h", test_cnt, test_data[test_cnt-1][31:0], r_data);
                    diff = 1;
                end
            end
            test_cnt <= test_cnt + 1;
        end
    end

    // 例化cache
    cache #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .WAY_NUM(WAY_NUM)
    ) cache_inst(
        .clk(clk),
        .rstn(rstn),
        .addr(addr),
        .r_req(r_req),
        .w_req(w_req),
        .w_data(w_data),
        .r_data(r_data),
        .miss(miss),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 内存
    mem #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH-LINE_OFFSET_WIDTH),
        .WAY_NUM(WAY_NUM)
    ) mem_inst(
        .clk(clk),
        .rstn(rstn),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 初始化测试数据
    initial begin
        test_addr[0] = 0;
        test_data[0] = 33'd7606690984;
        test_addr[1] = 32;
        test_data[1] = 33'd8035341310;
        test_addr[2] = 1;
        test_data[2] = 33'd1830337710;
        test_addr[3] = 2;
        test_data[3] = 33'd2722018698;
        test_addr[4] = 248;
        test_data[4] = 33'd995719055;
        test_addr[5] = 249;
        test_data[5] = 33'd3927970277;
        test_addr[6] = 250;
        test_data[6] = 33'd5697401980;
        test_addr[7] = 251;
        test_data[7] = 33'd5540123417;
        test_addr[8] = 3;
        test_data[8] = 33'd6390609751;
        test_addr[9] = 4;
        test_data[9] = 33'd340910773;
        test_addr[10] = 5;
        test_data[10] = 33'd426215752;
        test_addr[11] = 6;
        test_data[11] = 33'd7494251264;
        test_addr[12] = 7;
        test_data[12] = 33'd5261568043;
        test_addr[13] = 8;
        test_data[13] = 33'd8495106236;
        test_addr[14] = 9;
        test_data[14] = 33'd3430358658;
        test_addr[15] = 10;
        test_data[15] = 33'd6996403820;
        test_addr[16] = 11;
        test_data[16] = 33'd4437464051;
        test_addr[17] = 12;
        test_data[17] = 33'd1442523325;
        test_addr[18] = 13;
        test_data[18] = 33'd2440374455;
        test_addr[19] = 14;
        test_data[19] = 33'd1328303385;
        test_addr[20] = 15;
        test_data[20] = 33'd2428622533;
        test_addr[21] = 16;
        test_data[21] = 33'd38352283;
        test_addr[22] = 796;
        test_data[22] = 33'd4275211649;
        test_addr[23] = 17;
        test_data[23] = 33'd4627010622;
        test_addr[24] = 18;
        test_data[24] = 33'd5678085899;
        test_addr[25] = 19;
        test_data[25] = 33'd3066389384;
        test_addr[26] = 20;
        test_data[26] = 33'd6311232618;
        test_addr[27] = 21;
        test_data[27] = 33'd6299915841;
        test_addr[28] = 1019;
        test_data[28] = 33'd361342986;
        test_addr[29] = 22;
        test_data[29] = 33'd3991520861;
        test_addr[30] = 23;
        test_data[30] = 33'd4331393196;
        test_addr[31] = 24;
        test_data[31] = 33'd759408867;
        test_addr[32] = 25;
        test_data[32] = 33'd2632895408;
        test_addr[33] = 26;
        test_data[33] = 33'd3295931461;
        test_addr[34] = 27;
        test_data[34] = 33'd1081001156;
        test_addr[35] = 28;
        test_data[35] = 33'd1285008039;
        test_addr[36] = 613;
        test_data[36] = 33'd600314913;
        test_addr[37] = 614;
        test_data[37] = 33'd6401101506;
        test_addr[38] = 615;
        test_data[38] = 33'd4288664088;
        test_addr[39] = 616;
        test_data[39] = 33'd7345159614;
        test_addr[40] = 617;
        test_data[40] = 33'd6179479263;
        test_addr[41] = 618;
        test_data[41] = 33'd4559369986;
        test_addr[42] = 29;
        test_data[42] = 33'd943496892;
        test_addr[43] = 30;
        test_data[43] = 33'd7354103659;
        test_addr[44] = 31;
        test_data[44] = 33'd5470858984;
        test_addr[45] = 32;
        test_data[45] = 33'd3740374014;
        test_addr[46] = 33;
        test_data[46] = 33'd3213587532;
        test_addr[47] = 34;
        test_data[47] = 33'd3363095958;
        test_addr[48] = 35;
        test_data[48] = 33'd1763527796;
        test_addr[49] = 36;
        test_data[49] = 33'd6466514022;
        test_addr[50] = 37;
        test_data[50] = 33'd2923110415;
        test_addr[51] = 38;
        test_data[51] = 33'd8332460564;
        test_addr[52] = 39;
        test_data[52] = 33'd2019161959;
        test_addr[53] = 40;
        test_data[53] = 33'd8145729198;
        test_addr[54] = 41;
        test_data[54] = 33'd1144135439;
        test_addr[55] = 467;
        test_data[55] = 33'd1444845120;
        test_addr[56] = 468;
        test_data[56] = 33'd3544189000;
        test_addr[57] = 469;
        test_data[57] = 33'd821820080;
        test_addr[58] = 470;
        test_data[58] = 33'd5116981880;
        test_addr[59] = 471;
        test_data[59] = 33'd8393510425;
        test_addr[60] = 472;
        test_data[60] = 33'd1119598195;
        test_addr[61] = 473;
        test_data[61] = 33'd4114965494;
        test_addr[62] = 474;
        test_data[62] = 33'd2841812471;
        test_addr[63] = 475;
        test_data[63] = 33'd4470707941;
        test_addr[64] = 476;
        test_data[64] = 33'd1839489904;
        test_addr[65] = 477;
        test_data[65] = 33'd815049655;
        test_addr[66] = 478;
        test_data[66] = 33'd2289392119;
        test_addr[67] = 42;
        test_data[67] = 33'd7633741309;
        test_addr[68] = 43;
        test_data[68] = 33'd2969307118;
        test_addr[69] = 44;
        test_data[69] = 33'd3264450694;
        test_addr[70] = 45;
        test_data[70] = 33'd6929887853;
        test_addr[71] = 46;
        test_data[71] = 33'd7284918321;
        test_addr[72] = 47;
        test_data[72] = 33'd6571449605;
        test_addr[73] = 48;
        test_data[73] = 33'd3555854734;
        test_addr[74] = 440;
        test_data[74] = 33'd7501303376;
        test_addr[75] = 441;
        test_data[75] = 33'd6374578111;
        test_addr[76] = 442;
        test_data[76] = 33'd2950643337;
        test_addr[77] = 443;
        test_data[77] = 33'd1586603011;
        test_addr[78] = 49;
        test_data[78] = 33'd3795521150;
        test_addr[79] = 50;
        test_data[79] = 33'd3517050998;
        test_addr[80] = 290;
        test_data[80] = 33'd3645826661;
        test_addr[81] = 291;
        test_data[81] = 33'd2507289981;
        test_addr[82] = 292;
        test_data[82] = 33'd1640016259;
        test_addr[83] = 293;
        test_data[83] = 33'd1249044169;
        test_addr[84] = 294;
        test_data[84] = 33'd3223530803;
        test_addr[85] = 295;
        test_data[85] = 33'd1478684809;
        test_addr[86] = 296;
        test_data[86] = 33'd4661044283;
        test_addr[87] = 297;
        test_data[87] = 33'd2331663310;
        test_addr[88] = 298;
        test_data[88] = 33'd8475945775;
        test_addr[89] = 299;
        test_data[89] = 33'd2571156935;
        test_addr[90] = 300;
        test_data[90] = 33'd3281353580;
        test_addr[91] = 301;
        test_data[91] = 33'd4693308823;
        test_addr[92] = 51;
        test_data[92] = 33'd3196449230;
        test_addr[93] = 52;
        test_data[93] = 33'd1670309798;
        test_addr[94] = 53;
        test_data[94] = 33'd150061981;
        test_addr[95] = 748;
        test_data[95] = 33'd4371376208;
        test_addr[96] = 54;
        test_data[96] = 33'd586437743;
        test_addr[97] = 43;
        test_data[97] = 33'd6808980797;
        test_addr[98] = 55;
        test_data[98] = 33'd5897420755;
        test_addr[99] = 56;
        test_data[99] = 33'd4032767092;
        test_addr[100] = 57;
        test_data[100] = 33'd3015078990;
        test_addr[101] = 58;
        test_data[101] = 33'd2630100688;
        test_addr[102] = 59;
        test_data[102] = 33'd6854703267;
        test_addr[103] = 60;
        test_data[103] = 33'd6819120409;
        test_addr[104] = 61;
        test_data[104] = 33'd6874893096;
        test_addr[105] = 159;
        test_data[105] = 33'd3037698070;
        test_addr[106] = 160;
        test_data[106] = 33'd2288570994;
        test_addr[107] = 62;
        test_data[107] = 33'd304754323;
        test_addr[108] = 63;
        test_data[108] = 33'd1646915880;
        test_addr[109] = 64;
        test_data[109] = 33'd6261185364;
        test_addr[110] = 65;
        test_data[110] = 33'd1845517365;
        test_addr[111] = 66;
        test_data[111] = 33'd2814571527;
        test_addr[112] = 67;
        test_data[112] = 33'd7517214235;
        test_addr[113] = 68;
        test_data[113] = 33'd8364786480;
        test_addr[114] = 69;
        test_data[114] = 33'd5212554946;
        test_addr[115] = 70;
        test_data[115] = 33'd2049921272;
        test_addr[116] = 71;
        test_data[116] = 33'd2763155768;
        test_addr[117] = 72;
        test_data[117] = 33'd8208381171;
        test_addr[118] = 73;
        test_data[118] = 33'd404406686;
        test_addr[119] = 74;
        test_data[119] = 33'd3957199885;
        test_addr[120] = 593;
        test_data[120] = 33'd5365769197;
        test_addr[121] = 594;
        test_data[121] = 33'd7262593197;
        test_addr[122] = 595;
        test_data[122] = 33'd1646515767;
        test_addr[123] = 596;
        test_data[123] = 33'd2888243094;
        test_addr[124] = 597;
        test_data[124] = 33'd3535940700;
        test_addr[125] = 598;
        test_data[125] = 33'd5983850961;
        test_addr[126] = 599;
        test_data[126] = 33'd699313956;
        test_addr[127] = 600;
        test_data[127] = 33'd699365697;
        test_addr[128] = 601;
        test_data[128] = 33'd1061024359;
        test_addr[129] = 602;
        test_data[129] = 33'd523974119;
        test_addr[130] = 603;
        test_data[130] = 33'd1949152991;
        test_addr[131] = 604;
        test_data[131] = 33'd5408055643;
        test_addr[132] = 605;
        test_data[132] = 33'd1618144234;
        test_addr[133] = 606;
        test_data[133] = 33'd920782161;
        test_addr[134] = 607;
        test_data[134] = 33'd3986635328;
        test_addr[135] = 608;
        test_data[135] = 33'd2953791377;
        test_addr[136] = 609;
        test_data[136] = 33'd3511563354;
        test_addr[137] = 610;
        test_data[137] = 33'd2559326217;
        test_addr[138] = 611;
        test_data[138] = 33'd7236291049;
        test_addr[139] = 612;
        test_data[139] = 33'd702302819;
        test_addr[140] = 75;
        test_data[140] = 33'd869866033;
        test_addr[141] = 710;
        test_data[141] = 33'd5163249829;
        test_addr[142] = 711;
        test_data[142] = 33'd7409285638;
        test_addr[143] = 712;
        test_data[143] = 33'd265621438;
        test_addr[144] = 713;
        test_data[144] = 33'd3501601674;
        test_addr[145] = 714;
        test_data[145] = 33'd299549045;
        test_addr[146] = 715;
        test_data[146] = 33'd3297497505;
        test_addr[147] = 716;
        test_data[147] = 33'd292650974;
        test_addr[148] = 717;
        test_data[148] = 33'd4731578223;
        test_addr[149] = 718;
        test_data[149] = 33'd3656605274;
        test_addr[150] = 719;
        test_data[150] = 33'd602760059;
        test_addr[151] = 720;
        test_data[151] = 33'd264781874;
        test_addr[152] = 721;
        test_data[152] = 33'd4874270389;
        test_addr[153] = 722;
        test_data[153] = 33'd1583494039;
        test_addr[154] = 723;
        test_data[154] = 33'd7979458375;
        test_addr[155] = 724;
        test_data[155] = 33'd1061855659;
        test_addr[156] = 725;
        test_data[156] = 33'd5456939514;
        test_addr[157] = 726;
        test_data[157] = 33'd5775028576;
        test_addr[158] = 727;
        test_data[158] = 33'd2678040300;
        test_addr[159] = 728;
        test_data[159] = 33'd7117263844;
        test_addr[160] = 729;
        test_data[160] = 33'd4873753046;
        test_addr[161] = 730;
        test_data[161] = 33'd2998442618;
        test_addr[162] = 731;
        test_data[162] = 33'd3605685312;
        test_addr[163] = 732;
        test_data[163] = 33'd1766000469;
        test_addr[164] = 733;
        test_data[164] = 33'd3548136803;
        test_addr[165] = 734;
        test_data[165] = 33'd5606956066;
        test_addr[166] = 735;
        test_data[166] = 33'd8291843993;
        test_addr[167] = 736;
        test_data[167] = 33'd3833161201;
        test_addr[168] = 737;
        test_data[168] = 33'd7061190460;
        test_addr[169] = 738;
        test_data[169] = 33'd162191551;
        test_addr[170] = 76;
        test_data[170] = 33'd5378269558;
        test_addr[171] = 77;
        test_data[171] = 33'd2876543838;
        test_addr[172] = 78;
        test_data[172] = 33'd3671955214;
        test_addr[173] = 79;
        test_data[173] = 33'd238733017;
        test_addr[174] = 80;
        test_data[174] = 33'd2907114715;
        test_addr[175] = 81;
        test_data[175] = 33'd1759133022;
        test_addr[176] = 82;
        test_data[176] = 33'd2394041630;
        test_addr[177] = 83;
        test_data[177] = 33'd21120565;
        test_addr[178] = 84;
        test_data[178] = 33'd655204540;
        test_addr[179] = 85;
        test_data[179] = 33'd5982894112;
        test_addr[180] = 86;
        test_data[180] = 33'd88473128;
        test_addr[181] = 87;
        test_data[181] = 33'd5369349173;
        test_addr[182] = 88;
        test_data[182] = 33'd8440606319;
        test_addr[183] = 89;
        test_data[183] = 33'd227902140;
        test_addr[184] = 193;
        test_data[184] = 33'd1033777528;
        test_addr[185] = 194;
        test_data[185] = 33'd2955644450;
        test_addr[186] = 195;
        test_data[186] = 33'd6488813391;
        test_addr[187] = 196;
        test_data[187] = 33'd2584950764;
        test_addr[188] = 90;
        test_data[188] = 33'd7464669894;
        test_addr[189] = 91;
        test_data[189] = 33'd2419969866;
        test_addr[190] = 92;
        test_data[190] = 33'd6247480391;
        test_addr[191] = 93;
        test_data[191] = 33'd1228061459;
        test_addr[192] = 94;
        test_data[192] = 33'd3836173812;
        test_addr[193] = 95;
        test_data[193] = 33'd4605819778;
        test_addr[194] = 72;
        test_data[194] = 33'd5529516477;
        test_addr[195] = 73;
        test_data[195] = 33'd404406686;
        test_addr[196] = 96;
        test_data[196] = 33'd1615274362;
        test_addr[197] = 97;
        test_data[197] = 33'd3946323928;
        test_addr[198] = 98;
        test_data[198] = 33'd2576532341;
        test_addr[199] = 99;
        test_data[199] = 33'd3402368761;
        test_addr[200] = 100;
        test_data[200] = 33'd6329792614;
        test_addr[201] = 101;
        test_data[201] = 33'd4855307230;
        test_addr[202] = 102;
        test_data[202] = 33'd457023927;
        test_addr[203] = 103;
        test_data[203] = 33'd4732727241;
        test_addr[204] = 978;
        test_data[204] = 33'd2323391226;
        test_addr[205] = 979;
        test_data[205] = 33'd8255834368;
        test_addr[206] = 980;
        test_data[206] = 33'd3930060900;
        test_addr[207] = 981;
        test_data[207] = 33'd2623441966;
        test_addr[208] = 982;
        test_data[208] = 33'd6753596007;
        test_addr[209] = 983;
        test_data[209] = 33'd7955123158;
        test_addr[210] = 984;
        test_data[210] = 33'd5273898663;
        test_addr[211] = 985;
        test_data[211] = 33'd957211627;
        test_addr[212] = 986;
        test_data[212] = 33'd3822672388;
        test_addr[213] = 987;
        test_data[213] = 33'd1952340139;
        test_addr[214] = 988;
        test_data[214] = 33'd3995363066;
        test_addr[215] = 989;
        test_data[215] = 33'd4181739735;
        test_addr[216] = 990;
        test_data[216] = 33'd4853648795;
        test_addr[217] = 991;
        test_data[217] = 33'd88478458;
        test_addr[218] = 992;
        test_data[218] = 33'd669592020;
        test_addr[219] = 993;
        test_data[219] = 33'd1916779651;
        test_addr[220] = 104;
        test_data[220] = 33'd3745214105;
        test_addr[221] = 105;
        test_data[221] = 33'd3574643393;
        test_addr[222] = 106;
        test_data[222] = 33'd4071584875;
        test_addr[223] = 205;
        test_data[223] = 33'd4923192659;
        test_addr[224] = 206;
        test_data[224] = 33'd4213338333;
        test_addr[225] = 207;
        test_data[225] = 33'd513445133;
        test_addr[226] = 208;
        test_data[226] = 33'd3472524183;
        test_addr[227] = 107;
        test_data[227] = 33'd3862762663;
        test_addr[228] = 108;
        test_data[228] = 33'd2414169125;
        test_addr[229] = 109;
        test_data[229] = 33'd744992370;
        test_addr[230] = 110;
        test_data[230] = 33'd8177667470;
        test_addr[231] = 111;
        test_data[231] = 33'd1452439021;
        test_addr[232] = 112;
        test_data[232] = 33'd338946051;
        test_addr[233] = 113;
        test_data[233] = 33'd958838625;
        test_addr[234] = 114;
        test_data[234] = 33'd6673761826;
        test_addr[235] = 115;
        test_data[235] = 33'd1652892941;
        test_addr[236] = 28;
        test_data[236] = 33'd1285008039;
        test_addr[237] = 29;
        test_data[237] = 33'd943496892;
        test_addr[238] = 30;
        test_data[238] = 33'd3059136363;
        test_addr[239] = 31;
        test_data[239] = 33'd1175891688;
        test_addr[240] = 32;
        test_data[240] = 33'd3740374014;
        test_addr[241] = 33;
        test_data[241] = 33'd6812725625;
        test_addr[242] = 34;
        test_data[242] = 33'd3363095958;
        test_addr[243] = 35;
        test_data[243] = 33'd5509497068;
        test_addr[244] = 36;
        test_data[244] = 33'd6000069832;
        test_addr[245] = 37;
        test_data[245] = 33'd2923110415;
        test_addr[246] = 38;
        test_data[246] = 33'd4498804711;
        test_addr[247] = 39;
        test_data[247] = 33'd4377093961;
        test_addr[248] = 116;
        test_data[248] = 33'd3804836444;
        test_addr[249] = 117;
        test_data[249] = 33'd4220214550;
        test_addr[250] = 118;
        test_data[250] = 33'd5147239952;
        test_addr[251] = 119;
        test_data[251] = 33'd1527611154;
        test_addr[252] = 120;
        test_data[252] = 33'd2264552573;
        test_addr[253] = 121;
        test_data[253] = 33'd2605200182;
        test_addr[254] = 122;
        test_data[254] = 33'd3622924683;
        test_addr[255] = 123;
        test_data[255] = 33'd8510075084;
        test_addr[256] = 124;
        test_data[256] = 33'd4681634651;
        test_addr[257] = 125;
        test_data[257] = 33'd1528221139;
        test_addr[258] = 126;
        test_data[258] = 33'd4817449455;
        test_addr[259] = 127;
        test_data[259] = 33'd2531376941;
        test_addr[260] = 128;
        test_data[260] = 33'd4248669786;
        test_addr[261] = 129;
        test_data[261] = 33'd4507326927;
        test_addr[262] = 130;
        test_data[262] = 33'd3185392084;
        test_addr[263] = 131;
        test_data[263] = 33'd2412978687;
        test_addr[264] = 132;
        test_data[264] = 33'd347320602;
        test_addr[265] = 133;
        test_data[265] = 33'd5785944435;
        test_addr[266] = 134;
        test_data[266] = 33'd3657150815;
        test_addr[267] = 135;
        test_data[267] = 33'd1710980134;
        test_addr[268] = 136;
        test_data[268] = 33'd7646582444;
        test_addr[269] = 137;
        test_data[269] = 33'd3516062355;
        test_addr[270] = 138;
        test_data[270] = 33'd1254375529;
        test_addr[271] = 139;
        test_data[271] = 33'd8335175751;
        test_addr[272] = 140;
        test_data[272] = 33'd452007419;
        test_addr[273] = 141;
        test_data[273] = 33'd3732737218;
        test_addr[274] = 142;
        test_data[274] = 33'd5043358902;
        test_addr[275] = 143;
        test_data[275] = 33'd1991012920;
        test_addr[276] = 144;
        test_data[276] = 33'd6585631758;
        test_addr[277] = 145;
        test_data[277] = 33'd7250785548;
        test_addr[278] = 146;
        test_data[278] = 33'd2237304365;
        test_addr[279] = 147;
        test_data[279] = 33'd6203492183;
        test_addr[280] = 148;
        test_data[280] = 33'd7369101123;
        test_addr[281] = 149;
        test_data[281] = 33'd7097391914;
        test_addr[282] = 913;
        test_data[282] = 33'd2193415700;
        test_addr[283] = 914;
        test_data[283] = 33'd4579373040;
        test_addr[284] = 915;
        test_data[284] = 33'd5134752593;
        test_addr[285] = 916;
        test_data[285] = 33'd7414060854;
        test_addr[286] = 917;
        test_data[286] = 33'd2827507563;
        test_addr[287] = 918;
        test_data[287] = 33'd942389263;
        test_addr[288] = 919;
        test_data[288] = 33'd3709315097;
        test_addr[289] = 920;
        test_data[289] = 33'd7496566610;
        test_addr[290] = 150;
        test_data[290] = 33'd5864615448;
        test_addr[291] = 151;
        test_data[291] = 33'd5848900725;
        test_addr[292] = 152;
        test_data[292] = 33'd2253932096;
        test_addr[293] = 153;
        test_data[293] = 33'd3061874645;
        test_addr[294] = 154;
        test_data[294] = 33'd5833168323;
        test_addr[295] = 155;
        test_data[295] = 33'd1567660096;
        test_addr[296] = 156;
        test_data[296] = 33'd1564620619;
        test_addr[297] = 157;
        test_data[297] = 33'd2310668724;
        test_addr[298] = 158;
        test_data[298] = 33'd7851385812;
        test_addr[299] = 159;
        test_data[299] = 33'd3037698070;
        test_addr[300] = 160;
        test_data[300] = 33'd2288570994;
        test_addr[301] = 122;
        test_data[301] = 33'd3622924683;
        test_addr[302] = 123;
        test_data[302] = 33'd4215107788;
        test_addr[303] = 124;
        test_data[303] = 33'd386667355;
        test_addr[304] = 125;
        test_data[304] = 33'd5476970552;
        test_addr[305] = 126;
        test_data[305] = 33'd5284334937;
        test_addr[306] = 127;
        test_data[306] = 33'd6955723607;
        test_addr[307] = 128;
        test_data[307] = 33'd6411825664;
        test_addr[308] = 129;
        test_data[308] = 33'd212359631;
        test_addr[309] = 130;
        test_data[309] = 33'd3185392084;
        test_addr[310] = 131;
        test_data[310] = 33'd2412978687;
        test_addr[311] = 132;
        test_data[311] = 33'd4724981826;
        test_addr[312] = 133;
        test_data[312] = 33'd1490977139;
        test_addr[313] = 134;
        test_data[313] = 33'd3657150815;
        test_addr[314] = 135;
        test_data[314] = 33'd1710980134;
        test_addr[315] = 136;
        test_data[315] = 33'd3351615148;
        test_addr[316] = 137;
        test_data[316] = 33'd3516062355;
        test_addr[317] = 138;
        test_data[317] = 33'd1254375529;
        test_addr[318] = 139;
        test_data[318] = 33'd4040208455;
        test_addr[319] = 140;
        test_data[319] = 33'd452007419;
        test_addr[320] = 161;
        test_data[320] = 33'd2556436400;
        test_addr[321] = 162;
        test_data[321] = 33'd3143417896;
        test_addr[322] = 283;
        test_data[322] = 33'd2307617241;
        test_addr[323] = 284;
        test_data[323] = 33'd935136977;
        test_addr[324] = 285;
        test_data[324] = 33'd3139190243;
        test_addr[325] = 286;
        test_data[325] = 33'd2132904872;
        test_addr[326] = 287;
        test_data[326] = 33'd4288613521;
        test_addr[327] = 288;
        test_data[327] = 33'd2458363594;
        test_addr[328] = 289;
        test_data[328] = 33'd4124324693;
        test_addr[329] = 163;
        test_data[329] = 33'd3528470030;
        test_addr[330] = 164;
        test_data[330] = 33'd342696692;
        test_addr[331] = 165;
        test_data[331] = 33'd7892555770;
        test_addr[332] = 166;
        test_data[332] = 33'd2253906058;
        test_addr[333] = 167;
        test_data[333] = 33'd367704174;
        test_addr[334] = 168;
        test_data[334] = 33'd5159020181;
        test_addr[335] = 169;
        test_data[335] = 33'd705866065;
        test_addr[336] = 170;
        test_data[336] = 33'd911045719;
        test_addr[337] = 171;
        test_data[337] = 33'd4210643370;
        test_addr[338] = 172;
        test_data[338] = 33'd3645680872;
        test_addr[339] = 173;
        test_data[339] = 33'd1258215212;
        test_addr[340] = 174;
        test_data[340] = 33'd5447621970;
        test_addr[341] = 175;
        test_data[341] = 33'd3285653861;
        test_addr[342] = 176;
        test_data[342] = 33'd8201564937;
        test_addr[343] = 177;
        test_data[343] = 33'd6285953059;
        test_addr[344] = 178;
        test_data[344] = 33'd8173120189;
        test_addr[345] = 179;
        test_data[345] = 33'd487094244;
        test_addr[346] = 180;
        test_data[346] = 33'd1185846637;
        test_addr[347] = 181;
        test_data[347] = 33'd500375006;
        test_addr[348] = 182;
        test_data[348] = 33'd3172527317;
        test_addr[349] = 183;
        test_data[349] = 33'd5087909001;
        test_addr[350] = 184;
        test_data[350] = 33'd424689813;
        test_addr[351] = 185;
        test_data[351] = 33'd22147021;
        test_addr[352] = 763;
        test_data[352] = 33'd407903955;
        test_addr[353] = 764;
        test_data[353] = 33'd4591350789;
        test_addr[354] = 765;
        test_data[354] = 33'd6541836282;
        test_addr[355] = 766;
        test_data[355] = 33'd163370680;
        test_addr[356] = 767;
        test_data[356] = 33'd51594790;
        test_addr[357] = 768;
        test_data[357] = 33'd2995316459;
        test_addr[358] = 186;
        test_data[358] = 33'd3062031139;
        test_addr[359] = 187;
        test_data[359] = 33'd793217816;
        test_addr[360] = 188;
        test_data[360] = 33'd7577134065;
        test_addr[361] = 189;
        test_data[361] = 33'd669715075;
        test_addr[362] = 190;
        test_data[362] = 33'd1502392286;
        test_addr[363] = 191;
        test_data[363] = 33'd5518402837;
        test_addr[364] = 192;
        test_data[364] = 33'd4135019198;
        test_addr[365] = 193;
        test_data[365] = 33'd1033777528;
        test_addr[366] = 194;
        test_data[366] = 33'd2955644450;
        test_addr[367] = 195;
        test_data[367] = 33'd2193846095;
        test_addr[368] = 196;
        test_data[368] = 33'd2584950764;
        test_addr[369] = 197;
        test_data[369] = 33'd1696743885;
        test_addr[370] = 198;
        test_data[370] = 33'd2875093575;
        test_addr[371] = 199;
        test_data[371] = 33'd7572004240;
        test_addr[372] = 200;
        test_data[372] = 33'd8361762193;
        test_addr[373] = 201;
        test_data[373] = 33'd3316635280;
        test_addr[374] = 202;
        test_data[374] = 33'd5351836389;
        test_addr[375] = 203;
        test_data[375] = 33'd1831871360;
        test_addr[376] = 204;
        test_data[376] = 33'd1535612339;
        test_addr[377] = 205;
        test_data[377] = 33'd4677419096;
        test_addr[378] = 206;
        test_data[378] = 33'd4213338333;
        test_addr[379] = 207;
        test_data[379] = 33'd513445133;
        test_addr[380] = 208;
        test_data[380] = 33'd3472524183;
        test_addr[381] = 209;
        test_data[381] = 33'd7554045743;
        test_addr[382] = 210;
        test_data[382] = 33'd118596569;
        test_addr[383] = 211;
        test_data[383] = 33'd4202191155;
        test_addr[384] = 212;
        test_data[384] = 33'd2809482033;
        test_addr[385] = 213;
        test_data[385] = 33'd8143136555;
        test_addr[386] = 214;
        test_data[386] = 33'd635033231;
        test_addr[387] = 215;
        test_data[387] = 33'd4098659685;
        test_addr[388] = 216;
        test_data[388] = 33'd5876609870;
        test_addr[389] = 217;
        test_data[389] = 33'd2718828492;
        test_addr[390] = 218;
        test_data[390] = 33'd1056999408;
        test_addr[391] = 219;
        test_data[391] = 33'd193565387;
        test_addr[392] = 220;
        test_data[392] = 33'd6767738875;
        test_addr[393] = 221;
        test_data[393] = 33'd3019464660;
        test_addr[394] = 399;
        test_data[394] = 33'd509805444;
        test_addr[395] = 400;
        test_data[395] = 33'd6137275062;
        test_addr[396] = 401;
        test_data[396] = 33'd427139017;
        test_addr[397] = 402;
        test_data[397] = 33'd2447482056;
        test_addr[398] = 403;
        test_data[398] = 33'd5801213718;
        test_addr[399] = 404;
        test_data[399] = 33'd602052412;
        test_addr[400] = 405;
        test_data[400] = 33'd1195841942;
        test_addr[401] = 406;
        test_data[401] = 33'd532774694;
        test_addr[402] = 222;
        test_data[402] = 33'd1384897455;
        test_addr[403] = 223;
        test_data[403] = 33'd5676120780;
        test_addr[404] = 224;
        test_data[404] = 33'd463140193;
        test_addr[405] = 225;
        test_data[405] = 33'd5752618345;
        test_addr[406] = 226;
        test_data[406] = 33'd2717548623;
        test_addr[407] = 227;
        test_data[407] = 33'd2688484918;
        test_addr[408] = 228;
        test_data[408] = 33'd4120475529;
        test_addr[409] = 791;
        test_data[409] = 33'd1151411794;
        test_addr[410] = 792;
        test_data[410] = 33'd4897329810;
        test_addr[411] = 793;
        test_data[411] = 33'd8471763896;
        test_addr[412] = 794;
        test_data[412] = 33'd6155657428;
        test_addr[413] = 795;
        test_data[413] = 33'd2128607902;
        test_addr[414] = 796;
        test_data[414] = 33'd4275211649;
        test_addr[415] = 797;
        test_data[415] = 33'd115316762;
        test_addr[416] = 798;
        test_data[416] = 33'd4098353399;
        test_addr[417] = 799;
        test_data[417] = 33'd5813045251;
        test_addr[418] = 800;
        test_data[418] = 33'd754500382;
        test_addr[419] = 801;
        test_data[419] = 33'd3939763522;
        test_addr[420] = 802;
        test_data[420] = 33'd3959741461;
        test_addr[421] = 803;
        test_data[421] = 33'd2717076327;
        test_addr[422] = 804;
        test_data[422] = 33'd3891346024;
        test_addr[423] = 805;
        test_data[423] = 33'd571201105;
        test_addr[424] = 806;
        test_data[424] = 33'd5761441857;
        test_addr[425] = 807;
        test_data[425] = 33'd4934544759;
        test_addr[426] = 808;
        test_data[426] = 33'd158874295;
        test_addr[427] = 809;
        test_data[427] = 33'd8392787607;
        test_addr[428] = 810;
        test_data[428] = 33'd6275057515;
        test_addr[429] = 229;
        test_data[429] = 33'd665005425;
        test_addr[430] = 606;
        test_data[430] = 33'd920782161;
        test_addr[431] = 607;
        test_data[431] = 33'd3986635328;
        test_addr[432] = 608;
        test_data[432] = 33'd2953791377;
        test_addr[433] = 230;
        test_data[433] = 33'd5283425781;
        test_addr[434] = 231;
        test_data[434] = 33'd2346487764;
        test_addr[435] = 232;
        test_data[435] = 33'd6242430872;
        test_addr[436] = 233;
        test_data[436] = 33'd2492348860;
        test_addr[437] = 234;
        test_data[437] = 33'd3059098805;
        test_addr[438] = 235;
        test_data[438] = 33'd379016448;
        test_addr[439] = 236;
        test_data[439] = 33'd1954450839;
        test_addr[440] = 237;
        test_data[440] = 33'd3293190254;
        test_addr[441] = 238;
        test_data[441] = 33'd245166882;
        test_addr[442] = 239;
        test_data[442] = 33'd1677771600;
        test_addr[443] = 240;
        test_data[443] = 33'd524685732;
        test_addr[444] = 241;
        test_data[444] = 33'd3112036660;
        test_addr[445] = 242;
        test_data[445] = 33'd502196391;
        test_addr[446] = 243;
        test_data[446] = 33'd1440318250;
        test_addr[447] = 244;
        test_data[447] = 33'd1318439210;
        test_addr[448] = 245;
        test_data[448] = 33'd4619473625;
        test_addr[449] = 246;
        test_data[449] = 33'd801919684;
        test_addr[450] = 247;
        test_data[450] = 33'd3793934249;
        test_addr[451] = 248;
        test_data[451] = 33'd7367412845;
        test_addr[452] = 249;
        test_data[452] = 33'd7612050708;
        test_addr[453] = 250;
        test_data[453] = 33'd5882263129;
        test_addr[454] = 251;
        test_data[454] = 33'd1245156121;
        test_addr[455] = 252;
        test_data[455] = 33'd5149993689;
        test_addr[456] = 253;
        test_data[456] = 33'd2885822038;
        test_addr[457] = 254;
        test_data[457] = 33'd4395860666;
        test_addr[458] = 255;
        test_data[458] = 33'd3493356248;
        test_addr[459] = 256;
        test_data[459] = 33'd6839603523;
        test_addr[460] = 257;
        test_data[460] = 33'd3530939413;
        test_addr[461] = 436;
        test_data[461] = 33'd4034103201;
        test_addr[462] = 437;
        test_data[462] = 33'd465935354;
        test_addr[463] = 258;
        test_data[463] = 33'd1644063503;
        test_addr[464] = 873;
        test_data[464] = 33'd5425188702;
        test_addr[465] = 874;
        test_data[465] = 33'd5494589243;
        test_addr[466] = 875;
        test_data[466] = 33'd7212696707;
        test_addr[467] = 876;
        test_data[467] = 33'd3736677355;
        test_addr[468] = 877;
        test_data[468] = 33'd596443674;
        test_addr[469] = 878;
        test_data[469] = 33'd4315984434;
        test_addr[470] = 879;
        test_data[470] = 33'd4085858993;
        test_addr[471] = 880;
        test_data[471] = 33'd1009940429;
        test_addr[472] = 881;
        test_data[472] = 33'd3579846374;
        test_addr[473] = 882;
        test_data[473] = 33'd386405139;
        test_addr[474] = 883;
        test_data[474] = 33'd1933304197;
        test_addr[475] = 884;
        test_data[475] = 33'd6610350781;
        test_addr[476] = 259;
        test_data[476] = 33'd6628564951;
        test_addr[477] = 260;
        test_data[477] = 33'd1884041322;
        test_addr[478] = 261;
        test_data[478] = 33'd1776590124;
        test_addr[479] = 262;
        test_data[479] = 33'd7519644254;
        test_addr[480] = 263;
        test_data[480] = 33'd7495823252;
        test_addr[481] = 264;
        test_data[481] = 33'd4124826968;
        test_addr[482] = 265;
        test_data[482] = 33'd2848828629;
        test_addr[483] = 266;
        test_data[483] = 33'd2745001205;
        test_addr[484] = 267;
        test_data[484] = 33'd2501490696;
        test_addr[485] = 268;
        test_data[485] = 33'd4484051132;
        test_addr[486] = 269;
        test_data[486] = 33'd90054363;
        test_addr[487] = 270;
        test_data[487] = 33'd4155868294;
        test_addr[488] = 271;
        test_data[488] = 33'd1009868606;
        test_addr[489] = 272;
        test_data[489] = 33'd6627532733;
        test_addr[490] = 273;
        test_data[490] = 33'd3917527697;
        test_addr[491] = 274;
        test_data[491] = 33'd3059870078;
        test_addr[492] = 275;
        test_data[492] = 33'd5549593372;
        test_addr[493] = 276;
        test_data[493] = 33'd6763908993;
        test_addr[494] = 277;
        test_data[494] = 33'd5939450151;
        test_addr[495] = 278;
        test_data[495] = 33'd1532905441;
        test_addr[496] = 279;
        test_data[496] = 33'd8516134247;
        test_addr[497] = 280;
        test_data[497] = 33'd5219399924;
        test_addr[498] = 281;
        test_data[498] = 33'd3708121482;
        test_addr[499] = 282;
        test_data[499] = 33'd1881898418;
        test_addr[500] = 283;
        test_data[500] = 33'd2307617241;
        test_addr[501] = 284;
        test_data[501] = 33'd4900227638;
        test_addr[502] = 285;
        test_data[502] = 33'd3139190243;
        test_addr[503] = 286;
        test_data[503] = 33'd2132904872;
        test_addr[504] = 287;
        test_data[504] = 33'd4288613521;
        test_addr[505] = 288;
        test_data[505] = 33'd5194982214;
        test_addr[506] = 289;
        test_data[506] = 33'd4461592431;
        test_addr[507] = 290;
        test_data[507] = 33'd6333879931;
        test_addr[508] = 291;
        test_data[508] = 33'd2507289981;
        test_addr[509] = 292;
        test_data[509] = 33'd1640016259;
        test_addr[510] = 293;
        test_data[510] = 33'd1249044169;
        test_addr[511] = 294;
        test_data[511] = 33'd3223530803;
        test_addr[512] = 295;
        test_data[512] = 33'd1478684809;
        test_addr[513] = 296;
        test_data[513] = 33'd366076987;
        test_addr[514] = 297;
        test_data[514] = 33'd2331663310;
        test_addr[515] = 54;
        test_data[515] = 33'd586437743;
        test_addr[516] = 55;
        test_data[516] = 33'd7836776059;
        test_addr[517] = 298;
        test_data[517] = 33'd5019656995;
        test_addr[518] = 299;
        test_data[518] = 33'd2571156935;
        test_addr[519] = 300;
        test_data[519] = 33'd3281353580;
        test_addr[520] = 301;
        test_data[520] = 33'd7411472085;
        test_addr[521] = 302;
        test_data[521] = 33'd7952214281;
        test_addr[522] = 303;
        test_data[522] = 33'd4080236004;
        test_addr[523] = 304;
        test_data[523] = 33'd7915855285;
        test_addr[524] = 305;
        test_data[524] = 33'd405757788;
        test_addr[525] = 306;
        test_data[525] = 33'd3900608396;
        test_addr[526] = 307;
        test_data[526] = 33'd4032726540;
        test_addr[527] = 308;
        test_data[527] = 33'd4610159165;
        test_addr[528] = 309;
        test_data[528] = 33'd1432220972;
        test_addr[529] = 310;
        test_data[529] = 33'd727353973;
        test_addr[530] = 519;
        test_data[530] = 33'd8344465537;
        test_addr[531] = 520;
        test_data[531] = 33'd2563473161;
        test_addr[532] = 521;
        test_data[532] = 33'd3220870596;
        test_addr[533] = 522;
        test_data[533] = 33'd3048636483;
        test_addr[534] = 523;
        test_data[534] = 33'd2950126546;
        test_addr[535] = 524;
        test_data[535] = 33'd1326168490;
        test_addr[536] = 525;
        test_data[536] = 33'd6575983047;
        test_addr[537] = 526;
        test_data[537] = 33'd736640889;
        test_addr[538] = 527;
        test_data[538] = 33'd3884199812;
        test_addr[539] = 528;
        test_data[539] = 33'd7292332228;
        test_addr[540] = 529;
        test_data[540] = 33'd730554504;
        test_addr[541] = 530;
        test_data[541] = 33'd1157531596;
        test_addr[542] = 531;
        test_data[542] = 33'd6245766521;
        test_addr[543] = 532;
        test_data[543] = 33'd1996478713;
        test_addr[544] = 533;
        test_data[544] = 33'd1603575421;
        test_addr[545] = 534;
        test_data[545] = 33'd2544290285;
        test_addr[546] = 535;
        test_data[546] = 33'd1551618470;
        test_addr[547] = 536;
        test_data[547] = 33'd4216548472;
        test_addr[548] = 537;
        test_data[548] = 33'd1269482248;
        test_addr[549] = 538;
        test_data[549] = 33'd2662158238;
        test_addr[550] = 539;
        test_data[550] = 33'd1252831804;
        test_addr[551] = 540;
        test_data[551] = 33'd3769408227;
        test_addr[552] = 541;
        test_data[552] = 33'd3630666215;
        test_addr[553] = 542;
        test_data[553] = 33'd2523859335;
        test_addr[554] = 543;
        test_data[554] = 33'd108826463;
        test_addr[555] = 544;
        test_data[555] = 33'd8401130317;
        test_addr[556] = 545;
        test_data[556] = 33'd3521037345;
        test_addr[557] = 311;
        test_data[557] = 33'd261335557;
        test_addr[558] = 312;
        test_data[558] = 33'd2830282665;
        test_addr[559] = 313;
        test_data[559] = 33'd6753931465;
        test_addr[560] = 314;
        test_data[560] = 33'd303175971;
        test_addr[561] = 315;
        test_data[561] = 33'd735135208;
        test_addr[562] = 316;
        test_data[562] = 33'd4793188400;
        test_addr[563] = 317;
        test_data[563] = 33'd6669523364;
        test_addr[564] = 318;
        test_data[564] = 33'd2835077050;
        test_addr[565] = 465;
        test_data[565] = 33'd1435079633;
        test_addr[566] = 466;
        test_data[566] = 33'd2321964682;
        test_addr[567] = 319;
        test_data[567] = 33'd4652080533;
        test_addr[568] = 320;
        test_data[568] = 33'd2364460379;
        test_addr[569] = 747;
        test_data[569] = 33'd5282563425;
        test_addr[570] = 748;
        test_data[570] = 33'd76408912;
        test_addr[571] = 749;
        test_data[571] = 33'd821619415;
        test_addr[572] = 750;
        test_data[572] = 33'd1056728340;
        test_addr[573] = 321;
        test_data[573] = 33'd4756167202;
        test_addr[574] = 322;
        test_data[574] = 33'd2089037115;
        test_addr[575] = 305;
        test_data[575] = 33'd7591561464;
        test_addr[576] = 306;
        test_data[576] = 33'd3900608396;
        test_addr[577] = 307;
        test_data[577] = 33'd4439455076;
        test_addr[578] = 308;
        test_data[578] = 33'd315191869;
        test_addr[579] = 309;
        test_data[579] = 33'd6793077840;
        test_addr[580] = 310;
        test_data[580] = 33'd727353973;
        test_addr[581] = 311;
        test_data[581] = 33'd261335557;
        test_addr[582] = 312;
        test_data[582] = 33'd2830282665;
        test_addr[583] = 313;
        test_data[583] = 33'd2458964169;
        test_addr[584] = 314;
        test_data[584] = 33'd303175971;
        test_addr[585] = 315;
        test_data[585] = 33'd735135208;
        test_addr[586] = 316;
        test_data[586] = 33'd498221104;
        test_addr[587] = 317;
        test_data[587] = 33'd2374556068;
        test_addr[588] = 318;
        test_data[588] = 33'd2835077050;
        test_addr[589] = 319;
        test_data[589] = 33'd357113237;
        test_addr[590] = 320;
        test_data[590] = 33'd2364460379;
        test_addr[591] = 321;
        test_data[591] = 33'd461199906;
        test_addr[592] = 322;
        test_data[592] = 33'd4636303798;
        test_addr[593] = 323;
        test_data[593] = 33'd1861217836;
        test_addr[594] = 324;
        test_data[594] = 33'd7111776146;
        test_addr[595] = 325;
        test_data[595] = 33'd1715720789;
        test_addr[596] = 326;
        test_data[596] = 33'd3602797429;
        test_addr[597] = 327;
        test_data[597] = 33'd4382386232;
        test_addr[598] = 323;
        test_data[598] = 33'd1861217836;
        test_addr[599] = 324;
        test_data[599] = 33'd6252988741;
        test_addr[600] = 325;
        test_data[600] = 33'd6912582762;
        test_addr[601] = 326;
        test_data[601] = 33'd6982664022;
        test_addr[602] = 327;
        test_data[602] = 33'd5034294352;
        test_addr[603] = 328;
        test_data[603] = 33'd77460711;
        test_addr[604] = 329;
        test_data[604] = 33'd1741242015;
        test_addr[605] = 330;
        test_data[605] = 33'd3508612389;
        test_addr[606] = 331;
        test_data[606] = 33'd8524559031;
        test_addr[607] = 332;
        test_data[607] = 33'd4266769130;
        test_addr[608] = 786;
        test_data[608] = 33'd4292686456;
        test_addr[609] = 787;
        test_data[609] = 33'd6035210293;
        test_addr[610] = 788;
        test_data[610] = 33'd7434466733;
        test_addr[611] = 789;
        test_data[611] = 33'd1888095334;
        test_addr[612] = 790;
        test_data[612] = 33'd2157703382;
        test_addr[613] = 791;
        test_data[613] = 33'd1151411794;
        test_addr[614] = 792;
        test_data[614] = 33'd602362514;
        test_addr[615] = 793;
        test_data[615] = 33'd6577969704;
        test_addr[616] = 794;
        test_data[616] = 33'd7157612933;
        test_addr[617] = 795;
        test_data[617] = 33'd2128607902;
        test_addr[618] = 796;
        test_data[618] = 33'd4275211649;
        test_addr[619] = 797;
        test_data[619] = 33'd7857155032;
        test_addr[620] = 798;
        test_data[620] = 33'd4098353399;
        test_addr[621] = 799;
        test_data[621] = 33'd1518077955;
        test_addr[622] = 800;
        test_data[622] = 33'd754500382;
        test_addr[623] = 801;
        test_data[623] = 33'd4879361151;
        test_addr[624] = 802;
        test_data[624] = 33'd7358192512;
        test_addr[625] = 803;
        test_data[625] = 33'd5329739779;
        test_addr[626] = 804;
        test_data[626] = 33'd7780273057;
        test_addr[627] = 805;
        test_data[627] = 33'd6813106752;
        test_addr[628] = 806;
        test_data[628] = 33'd1466474561;
        test_addr[629] = 807;
        test_data[629] = 33'd639577463;
        test_addr[630] = 808;
        test_data[630] = 33'd158874295;
        test_addr[631] = 809;
        test_data[631] = 33'd8263297119;
        test_addr[632] = 810;
        test_data[632] = 33'd1980090219;
        test_addr[633] = 811;
        test_data[633] = 33'd7263779840;
        test_addr[634] = 812;
        test_data[634] = 33'd1965390572;
        test_addr[635] = 813;
        test_data[635] = 33'd7502366644;
        test_addr[636] = 814;
        test_data[636] = 33'd2532614522;
        test_addr[637] = 815;
        test_data[637] = 33'd116081840;
        test_addr[638] = 816;
        test_data[638] = 33'd2089907260;
        test_addr[639] = 817;
        test_data[639] = 33'd6622016559;
        test_addr[640] = 818;
        test_data[640] = 33'd1746275809;
        test_addr[641] = 819;
        test_data[641] = 33'd7702299705;
        test_addr[642] = 820;
        test_data[642] = 33'd3200758228;
        test_addr[643] = 821;
        test_data[643] = 33'd4426857976;
        test_addr[644] = 822;
        test_data[644] = 33'd2790105153;
        test_addr[645] = 823;
        test_data[645] = 33'd2118102746;
        test_addr[646] = 824;
        test_data[646] = 33'd4185437212;
        test_addr[647] = 825;
        test_data[647] = 33'd1444494147;
        test_addr[648] = 826;
        test_data[648] = 33'd4957417803;
        test_addr[649] = 827;
        test_data[649] = 33'd4271161680;
        test_addr[650] = 828;
        test_data[650] = 33'd3143336390;
        test_addr[651] = 829;
        test_data[651] = 33'd2471067861;
        test_addr[652] = 830;
        test_data[652] = 33'd2151514164;
        test_addr[653] = 831;
        test_data[653] = 33'd3512387836;
        test_addr[654] = 832;
        test_data[654] = 33'd2442866266;
        test_addr[655] = 833;
        test_data[655] = 33'd807590553;
        test_addr[656] = 333;
        test_data[656] = 33'd2296982685;
        test_addr[657] = 334;
        test_data[657] = 33'd2783766917;
        test_addr[658] = 335;
        test_data[658] = 33'd1195626943;
        test_addr[659] = 336;
        test_data[659] = 33'd1688024943;
        test_addr[660] = 337;
        test_data[660] = 33'd5045228725;
        test_addr[661] = 338;
        test_data[661] = 33'd1821314294;
        test_addr[662] = 339;
        test_data[662] = 33'd3023854751;
        test_addr[663] = 340;
        test_data[663] = 33'd1638179589;
        test_addr[664] = 341;
        test_data[664] = 33'd315843574;
        test_addr[665] = 342;
        test_data[665] = 33'd4363622697;
        test_addr[666] = 343;
        test_data[666] = 33'd2846218665;
        test_addr[667] = 344;
        test_data[667] = 33'd5063190739;
        test_addr[668] = 345;
        test_data[668] = 33'd2791959723;
        test_addr[669] = 346;
        test_data[669] = 33'd3770003965;
        test_addr[670] = 35;
        test_data[670] = 33'd1214529772;
        test_addr[671] = 36;
        test_data[671] = 33'd1705102536;
        test_addr[672] = 37;
        test_data[672] = 33'd8187440079;
        test_addr[673] = 38;
        test_data[673] = 33'd203837415;
        test_addr[674] = 39;
        test_data[674] = 33'd6014591401;
        test_addr[675] = 40;
        test_data[675] = 33'd4472815509;
        test_addr[676] = 41;
        test_data[676] = 33'd1144135439;
        test_addr[677] = 42;
        test_data[677] = 33'd5169766887;
        test_addr[678] = 43;
        test_data[678] = 33'd2514013501;
        test_addr[679] = 44;
        test_data[679] = 33'd3264450694;
        test_addr[680] = 45;
        test_data[680] = 33'd4419299524;
        test_addr[681] = 46;
        test_data[681] = 33'd2989951025;
        test_addr[682] = 47;
        test_data[682] = 33'd2276482309;
        test_addr[683] = 48;
        test_data[683] = 33'd8132577458;
        test_addr[684] = 49;
        test_data[684] = 33'd3795521150;
        test_addr[685] = 50;
        test_data[685] = 33'd3517050998;
        test_addr[686] = 51;
        test_data[686] = 33'd8260922654;
        test_addr[687] = 52;
        test_data[687] = 33'd1670309798;
        test_addr[688] = 53;
        test_data[688] = 33'd5449431887;
        test_addr[689] = 347;
        test_data[689] = 33'd4150740891;
        test_addr[690] = 348;
        test_data[690] = 33'd904943400;
        test_addr[691] = 349;
        test_data[691] = 33'd3103175904;
        test_addr[692] = 350;
        test_data[692] = 33'd4912190208;
        test_addr[693] = 351;
        test_data[693] = 33'd2365388450;
        test_addr[694] = 352;
        test_data[694] = 33'd163922335;
        test_addr[695] = 353;
        test_data[695] = 33'd3565100911;
        test_addr[696] = 354;
        test_data[696] = 33'd8375945166;
        test_addr[697] = 355;
        test_data[697] = 33'd3917761171;
        test_addr[698] = 356;
        test_data[698] = 33'd2257235136;
        test_addr[699] = 357;
        test_data[699] = 33'd3927443995;
        test_addr[700] = 358;
        test_data[700] = 33'd3685422029;
        test_addr[701] = 359;
        test_data[701] = 33'd3154057553;
        test_addr[702] = 360;
        test_data[702] = 33'd3069921140;
        test_addr[703] = 361;
        test_data[703] = 33'd5694896564;
        test_addr[704] = 362;
        test_data[704] = 33'd2935077560;
        test_addr[705] = 363;
        test_data[705] = 33'd2723076636;
        test_addr[706] = 364;
        test_data[706] = 33'd1333182938;
        test_addr[707] = 365;
        test_data[707] = 33'd1161783265;
        test_addr[708] = 366;
        test_data[708] = 33'd7294106957;
        test_addr[709] = 367;
        test_data[709] = 33'd1351470440;
        test_addr[710] = 368;
        test_data[710] = 33'd4078620521;
        test_addr[711] = 369;
        test_data[711] = 33'd6402962279;
        test_addr[712] = 370;
        test_data[712] = 33'd4446799408;
        test_addr[713] = 371;
        test_data[713] = 33'd2775974076;
        test_addr[714] = 372;
        test_data[714] = 33'd3653485486;
        test_addr[715] = 373;
        test_data[715] = 33'd3628187523;
        test_addr[716] = 374;
        test_data[716] = 33'd8377038502;
        test_addr[717] = 375;
        test_data[717] = 33'd2719622023;
        test_addr[718] = 376;
        test_data[718] = 33'd6560213559;
        test_addr[719] = 377;
        test_data[719] = 33'd436835430;
        test_addr[720] = 378;
        test_data[720] = 33'd515798227;
        test_addr[721] = 379;
        test_data[721] = 33'd708784957;
        test_addr[722] = 380;
        test_data[722] = 33'd1150466899;
        test_addr[723] = 381;
        test_data[723] = 33'd1741094807;
        test_addr[724] = 382;
        test_data[724] = 33'd3223401649;
        test_addr[725] = 383;
        test_data[725] = 33'd5379240956;
        test_addr[726] = 384;
        test_data[726] = 33'd4847637602;
        test_addr[727] = 385;
        test_data[727] = 33'd817202464;
        test_addr[728] = 402;
        test_data[728] = 33'd2447482056;
        test_addr[729] = 403;
        test_data[729] = 33'd1506246422;
        test_addr[730] = 404;
        test_data[730] = 33'd4423927561;
        test_addr[731] = 405;
        test_data[731] = 33'd6248911872;
        test_addr[732] = 406;
        test_data[732] = 33'd532774694;
        test_addr[733] = 386;
        test_data[733] = 33'd1481982667;
        test_addr[734] = 387;
        test_data[734] = 33'd5886239441;
        test_addr[735] = 388;
        test_data[735] = 33'd3781905541;
        test_addr[736] = 389;
        test_data[736] = 33'd3497432784;
        test_addr[737] = 390;
        test_data[737] = 33'd5757528485;
        test_addr[738] = 391;
        test_data[738] = 33'd3183432554;
        test_addr[739] = 392;
        test_data[739] = 33'd2117412331;
        test_addr[740] = 357;
        test_data[740] = 33'd3927443995;
        test_addr[741] = 358;
        test_data[741] = 33'd3685422029;
        test_addr[742] = 359;
        test_data[742] = 33'd3154057553;
        test_addr[743] = 360;
        test_data[743] = 33'd3069921140;
        test_addr[744] = 361;
        test_data[744] = 33'd6709518393;
        test_addr[745] = 362;
        test_data[745] = 33'd7368239602;
        test_addr[746] = 363;
        test_data[746] = 33'd2723076636;
        test_addr[747] = 364;
        test_data[747] = 33'd1333182938;
        test_addr[748] = 365;
        test_data[748] = 33'd1161783265;
        test_addr[749] = 366;
        test_data[749] = 33'd2999139661;
        test_addr[750] = 367;
        test_data[750] = 33'd7721450560;
        test_addr[751] = 368;
        test_data[751] = 33'd4679368881;
        test_addr[752] = 369;
        test_data[752] = 33'd2107994983;
        test_addr[753] = 370;
        test_data[753] = 33'd151832112;
        test_addr[754] = 371;
        test_data[754] = 33'd2775974076;
        test_addr[755] = 372;
        test_data[755] = 33'd3653485486;
        test_addr[756] = 373;
        test_data[756] = 33'd6011706928;
        test_addr[757] = 374;
        test_data[757] = 33'd4082071206;
        test_addr[758] = 393;
        test_data[758] = 33'd479449245;
        test_addr[759] = 394;
        test_data[759] = 33'd4514910212;
        test_addr[760] = 395;
        test_data[760] = 33'd7974474962;
        test_addr[761] = 396;
        test_data[761] = 33'd4418666684;
        test_addr[762] = 397;
        test_data[762] = 33'd8435965737;
        test_addr[763] = 398;
        test_data[763] = 33'd3505084960;
        test_addr[764] = 399;
        test_data[764] = 33'd5539813442;
        test_addr[765] = 400;
        test_data[765] = 33'd7778887110;
        test_addr[766] = 401;
        test_data[766] = 33'd427139017;
        test_addr[767] = 402;
        test_data[767] = 33'd5498352345;
        test_addr[768] = 403;
        test_data[768] = 33'd4829720894;
        test_addr[769] = 404;
        test_data[769] = 33'd128960265;
        test_addr[770] = 405;
        test_data[770] = 33'd5181447959;
        test_addr[771] = 406;
        test_data[771] = 33'd5694739807;
        test_addr[772] = 407;
        test_data[772] = 33'd7945948717;
        test_addr[773] = 408;
        test_data[773] = 33'd1991242564;
        test_addr[774] = 409;
        test_data[774] = 33'd881702054;
        test_addr[775] = 142;
        test_data[775] = 33'd7173355747;
        test_addr[776] = 143;
        test_data[776] = 33'd4302682330;
        test_addr[777] = 144;
        test_data[777] = 33'd5660486463;
        test_addr[778] = 145;
        test_data[778] = 33'd2955818252;
        test_addr[779] = 146;
        test_data[779] = 33'd4406178750;
        test_addr[780] = 410;
        test_data[780] = 33'd3442998655;
        test_addr[781] = 411;
        test_data[781] = 33'd2509072348;
        test_addr[782] = 412;
        test_data[782] = 33'd3063633923;
        test_addr[783] = 413;
        test_data[783] = 33'd4263007220;
        test_addr[784] = 414;
        test_data[784] = 33'd2622463751;
        test_addr[785] = 415;
        test_data[785] = 33'd2483981373;
        test_addr[786] = 416;
        test_data[786] = 33'd3762483973;
        test_addr[787] = 417;
        test_data[787] = 33'd857483597;
        test_addr[788] = 418;
        test_data[788] = 33'd3304050455;
        test_addr[789] = 419;
        test_data[789] = 33'd3868382538;
        test_addr[790] = 420;
        test_data[790] = 33'd2008269494;
        test_addr[791] = 421;
        test_data[791] = 33'd3124744987;
        test_addr[792] = 422;
        test_data[792] = 33'd2139306794;
        test_addr[793] = 423;
        test_data[793] = 33'd7396574049;
        test_addr[794] = 424;
        test_data[794] = 33'd4107482093;
        test_addr[795] = 425;
        test_data[795] = 33'd6741685948;
        test_addr[796] = 426;
        test_data[796] = 33'd7391331744;
        test_addr[797] = 427;
        test_data[797] = 33'd1334217002;
        test_addr[798] = 428;
        test_data[798] = 33'd807619004;
        test_addr[799] = 429;
        test_data[799] = 33'd8389601540;
        test_addr[800] = 430;
        test_data[800] = 33'd896214945;
        test_addr[801] = 431;
        test_data[801] = 33'd3279784998;
        test_addr[802] = 432;
        test_data[802] = 33'd842198295;
        test_addr[803] = 433;
        test_data[803] = 33'd5824821207;
        test_addr[804] = 434;
        test_data[804] = 33'd4717968449;
        test_addr[805] = 562;
        test_data[805] = 33'd3011983409;
        test_addr[806] = 563;
        test_data[806] = 33'd3434699751;
        test_addr[807] = 564;
        test_data[807] = 33'd869541130;
        test_addr[808] = 565;
        test_data[808] = 33'd1601476386;
        test_addr[809] = 566;
        test_data[809] = 33'd6847110926;
        test_addr[810] = 567;
        test_data[810] = 33'd8271247447;
        test_addr[811] = 435;
        test_data[811] = 33'd2315575124;
        test_addr[812] = 436;
        test_data[812] = 33'd4034103201;
        test_addr[813] = 437;
        test_data[813] = 33'd6598093794;
        test_addr[814] = 438;
        test_data[814] = 33'd636048466;
        test_addr[815] = 439;
        test_data[815] = 33'd7482274907;
        test_addr[816] = 440;
        test_data[816] = 33'd5026354572;
        test_addr[817] = 441;
        test_data[817] = 33'd2079610815;
        test_addr[818] = 442;
        test_data[818] = 33'd2950643337;
        test_addr[819] = 443;
        test_data[819] = 33'd1586603011;
        test_addr[820] = 444;
        test_data[820] = 33'd2677223067;
        test_addr[821] = 445;
        test_data[821] = 33'd4932013754;
        test_addr[822] = 446;
        test_data[822] = 33'd1320511667;
        test_addr[823] = 447;
        test_data[823] = 33'd3084548448;
        test_addr[824] = 448;
        test_data[824] = 33'd2047532963;
        test_addr[825] = 449;
        test_data[825] = 33'd658651725;
        test_addr[826] = 450;
        test_data[826] = 33'd2853006304;
        test_addr[827] = 451;
        test_data[827] = 33'd5067342673;
        test_addr[828] = 452;
        test_data[828] = 33'd1012981055;
        test_addr[829] = 453;
        test_data[829] = 33'd4144249236;
        test_addr[830] = 565;
        test_data[830] = 33'd1601476386;
        test_addr[831] = 566;
        test_data[831] = 33'd2552143630;
        test_addr[832] = 567;
        test_data[832] = 33'd3976280151;
        test_addr[833] = 568;
        test_data[833] = 33'd1475611248;
        test_addr[834] = 569;
        test_data[834] = 33'd4859379060;
        test_addr[835] = 570;
        test_data[835] = 33'd4180903970;
        test_addr[836] = 571;
        test_data[836] = 33'd8143447028;
        test_addr[837] = 572;
        test_data[837] = 33'd403146832;
        test_addr[838] = 573;
        test_data[838] = 33'd660266423;
        test_addr[839] = 454;
        test_data[839] = 33'd7301450849;
        test_addr[840] = 455;
        test_data[840] = 33'd4791580;
        test_addr[841] = 456;
        test_data[841] = 33'd2010861474;
        test_addr[842] = 457;
        test_data[842] = 33'd4310737026;
        test_addr[843] = 33;
        test_data[843] = 33'd6303559338;
        test_addr[844] = 34;
        test_data[844] = 33'd3363095958;
        test_addr[845] = 35;
        test_data[845] = 33'd4770688275;
        test_addr[846] = 36;
        test_data[846] = 33'd8307190261;
        test_addr[847] = 37;
        test_data[847] = 33'd7650091424;
        test_addr[848] = 38;
        test_data[848] = 33'd203837415;
        test_addr[849] = 39;
        test_data[849] = 33'd5759794428;
        test_addr[850] = 40;
        test_data[850] = 33'd177848213;
        test_addr[851] = 41;
        test_data[851] = 33'd1144135439;
        test_addr[852] = 42;
        test_data[852] = 33'd7979377105;
        test_addr[853] = 43;
        test_data[853] = 33'd2514013501;
        test_addr[854] = 44;
        test_data[854] = 33'd3264450694;
        test_addr[855] = 45;
        test_data[855] = 33'd124332228;
        test_addr[856] = 46;
        test_data[856] = 33'd5028885415;
        test_addr[857] = 47;
        test_data[857] = 33'd2276482309;
        test_addr[858] = 48;
        test_data[858] = 33'd3837610162;
        test_addr[859] = 49;
        test_data[859] = 33'd3795521150;
        test_addr[860] = 50;
        test_data[860] = 33'd3517050998;
        test_addr[861] = 51;
        test_data[861] = 33'd3965955358;
        test_addr[862] = 52;
        test_data[862] = 33'd1670309798;
        test_addr[863] = 53;
        test_data[863] = 33'd6054698775;
        test_addr[864] = 54;
        test_data[864] = 33'd8057163735;
        test_addr[865] = 458;
        test_data[865] = 33'd4143306261;
        test_addr[866] = 459;
        test_data[866] = 33'd1894780540;
        test_addr[867] = 460;
        test_data[867] = 33'd7010493793;
        test_addr[868] = 461;
        test_data[868] = 33'd6502477574;
        test_addr[869] = 462;
        test_data[869] = 33'd2318869365;
        test_addr[870] = 463;
        test_data[870] = 33'd909928079;
        test_addr[871] = 38;
        test_data[871] = 33'd203837415;
        test_addr[872] = 464;
        test_data[872] = 33'd3521762258;
        test_addr[873] = 465;
        test_data[873] = 33'd8468289526;
        test_addr[874] = 466;
        test_data[874] = 33'd5886584618;
        test_addr[875] = 467;
        test_data[875] = 33'd1444845120;
        test_addr[876] = 85;
        test_data[876] = 33'd8403486630;
        test_addr[877] = 86;
        test_data[877] = 33'd5200228362;
        test_addr[878] = 87;
        test_data[878] = 33'd1074381877;
        test_addr[879] = 88;
        test_data[879] = 33'd4145639023;
        test_addr[880] = 89;
        test_data[880] = 33'd7697268760;
        test_addr[881] = 90;
        test_data[881] = 33'd3169702598;
        test_addr[882] = 91;
        test_data[882] = 33'd2419969866;
        test_addr[883] = 468;
        test_data[883] = 33'd3544189000;
        test_addr[884] = 469;
        test_data[884] = 33'd821820080;
        test_addr[885] = 470;
        test_data[885] = 33'd822014584;
        test_addr[886] = 471;
        test_data[886] = 33'd4098543129;
        test_addr[887] = 472;
        test_data[887] = 33'd6441422387;
        test_addr[888] = 473;
        test_data[888] = 33'd4114965494;
        test_addr[889] = 474;
        test_data[889] = 33'd2841812471;
        test_addr[890] = 475;
        test_data[890] = 33'd175740645;
        test_addr[891] = 385;
        test_data[891] = 33'd817202464;
        test_addr[892] = 386;
        test_data[892] = 33'd7336373828;
        test_addr[893] = 387;
        test_data[893] = 33'd1591272145;
        test_addr[894] = 388;
        test_data[894] = 33'd3781905541;
        test_addr[895] = 389;
        test_data[895] = 33'd3497432784;
        test_addr[896] = 390;
        test_data[896] = 33'd6838727960;
        test_addr[897] = 391;
        test_data[897] = 33'd4484725021;
        test_addr[898] = 392;
        test_data[898] = 33'd5301651977;
        test_addr[899] = 476;
        test_data[899] = 33'd1839489904;
        test_addr[900] = 477;
        test_data[900] = 33'd815049655;
        test_addr[901] = 478;
        test_data[901] = 33'd2289392119;
        test_addr[902] = 479;
        test_data[902] = 33'd6359983561;
        test_addr[903] = 480;
        test_data[903] = 33'd125390000;
        test_addr[904] = 481;
        test_data[904] = 33'd2639408353;
        test_addr[905] = 482;
        test_data[905] = 33'd3393357937;
        test_addr[906] = 483;
        test_data[906] = 33'd5618092133;
        test_addr[907] = 484;
        test_data[907] = 33'd998179708;
        test_addr[908] = 184;
        test_data[908] = 33'd424689813;
        test_addr[909] = 185;
        test_data[909] = 33'd6686366701;
        test_addr[910] = 186;
        test_data[910] = 33'd3062031139;
        test_addr[911] = 187;
        test_data[911] = 33'd793217816;
        test_addr[912] = 188;
        test_data[912] = 33'd4987152450;
        test_addr[913] = 189;
        test_data[913] = 33'd7036357792;
        test_addr[914] = 190;
        test_data[914] = 33'd7969514703;
        test_addr[915] = 191;
        test_data[915] = 33'd1223435541;
        test_addr[916] = 192;
        test_data[916] = 33'd4986412806;
        test_addr[917] = 193;
        test_data[917] = 33'd1033777528;
        test_addr[918] = 194;
        test_data[918] = 33'd2955644450;
        test_addr[919] = 195;
        test_data[919] = 33'd2193846095;
        test_addr[920] = 196;
        test_data[920] = 33'd2584950764;
        test_addr[921] = 197;
        test_data[921] = 33'd1696743885;
        test_addr[922] = 198;
        test_data[922] = 33'd2875093575;
        test_addr[923] = 199;
        test_data[923] = 33'd4412835605;
        test_addr[924] = 200;
        test_data[924] = 33'd4066794897;
        test_addr[925] = 201;
        test_data[925] = 33'd3316635280;
        test_addr[926] = 202;
        test_data[926] = 33'd1056869093;
        test_addr[927] = 203;
        test_data[927] = 33'd1831871360;
        test_addr[928] = 204;
        test_data[928] = 33'd7172758867;
        test_addr[929] = 205;
        test_data[929] = 33'd382451800;
        test_addr[930] = 206;
        test_data[930] = 33'd4213338333;
        test_addr[931] = 207;
        test_data[931] = 33'd513445133;
        test_addr[932] = 208;
        test_data[932] = 33'd3472524183;
        test_addr[933] = 485;
        test_data[933] = 33'd1497784997;
        test_addr[934] = 486;
        test_data[934] = 33'd3551446877;
        test_addr[935] = 774;
        test_data[935] = 33'd3061105897;
        test_addr[936] = 487;
        test_data[936] = 33'd8528891704;
        test_addr[937] = 488;
        test_data[937] = 33'd3230286556;
        test_addr[938] = 489;
        test_data[938] = 33'd654573334;
        test_addr[939] = 490;
        test_data[939] = 33'd4090258182;
        test_addr[940] = 491;
        test_data[940] = 33'd2199790567;
        test_addr[941] = 492;
        test_data[941] = 33'd2583156540;
        test_addr[942] = 493;
        test_data[942] = 33'd2115438628;
        test_addr[943] = 494;
        test_data[943] = 33'd4244092772;
        test_addr[944] = 495;
        test_data[944] = 33'd4312288548;
        test_addr[945] = 496;
        test_data[945] = 33'd7332507496;
        test_addr[946] = 497;
        test_data[946] = 33'd3663618438;
        test_addr[947] = 489;
        test_data[947] = 33'd654573334;
        test_addr[948] = 498;
        test_data[948] = 33'd4163492510;
        test_addr[949] = 499;
        test_data[949] = 33'd5351167369;
        test_addr[950] = 500;
        test_data[950] = 33'd5815338621;
        test_addr[951] = 501;
        test_data[951] = 33'd2592532499;
        test_addr[952] = 502;
        test_data[952] = 33'd1661402023;
        test_addr[953] = 503;
        test_data[953] = 33'd1431025879;
        test_addr[954] = 504;
        test_data[954] = 33'd225331988;
        test_addr[955] = 505;
        test_data[955] = 33'd5272953874;
        test_addr[956] = 506;
        test_data[956] = 33'd7773975940;
        test_addr[957] = 507;
        test_data[957] = 33'd3984605869;
        test_addr[958] = 508;
        test_data[958] = 33'd1247575968;
        test_addr[959] = 509;
        test_data[959] = 33'd1995849586;
        test_addr[960] = 510;
        test_data[960] = 33'd513403764;
        test_addr[961] = 511;
        test_data[961] = 33'd4030006546;
        test_addr[962] = 512;
        test_data[962] = 33'd1581423827;
        test_addr[963] = 513;
        test_data[963] = 33'd421452164;
        test_addr[964] = 514;
        test_data[964] = 33'd2973446334;
        test_addr[965] = 515;
        test_data[965] = 33'd4209937496;
        test_addr[966] = 516;
        test_data[966] = 33'd1918061132;
        test_addr[967] = 517;
        test_data[967] = 33'd4067077614;
        test_addr[968] = 518;
        test_data[968] = 33'd849664853;
        test_addr[969] = 519;
        test_data[969] = 33'd4049498241;
        test_addr[970] = 520;
        test_data[970] = 33'd7520293385;
        test_addr[971] = 521;
        test_data[971] = 33'd3220870596;
        test_addr[972] = 522;
        test_data[972] = 33'd3048636483;
        test_addr[973] = 523;
        test_data[973] = 33'd5677818763;
        test_addr[974] = 524;
        test_data[974] = 33'd4870462325;
        test_addr[975] = 525;
        test_data[975] = 33'd2281015751;
        test_addr[976] = 526;
        test_data[976] = 33'd736640889;
        test_addr[977] = 636;
        test_data[977] = 33'd6259078961;
        test_addr[978] = 637;
        test_data[978] = 33'd7437032199;
        test_addr[979] = 638;
        test_data[979] = 33'd3568991821;
        test_addr[980] = 639;
        test_data[980] = 33'd8357145113;
        test_addr[981] = 640;
        test_data[981] = 33'd3889086438;
        test_addr[982] = 641;
        test_data[982] = 33'd3812820741;
        test_addr[983] = 642;
        test_data[983] = 33'd5277207304;
        test_addr[984] = 643;
        test_data[984] = 33'd6535139394;
        test_addr[985] = 644;
        test_data[985] = 33'd7324355419;
        test_addr[986] = 645;
        test_data[986] = 33'd4494856756;
        test_addr[987] = 646;
        test_data[987] = 33'd5620256829;
        test_addr[988] = 647;
        test_data[988] = 33'd5598409569;
        test_addr[989] = 648;
        test_data[989] = 33'd2300180881;
        test_addr[990] = 649;
        test_data[990] = 33'd8542392617;
        test_addr[991] = 650;
        test_data[991] = 33'd2784853932;
        test_addr[992] = 651;
        test_data[992] = 33'd7683143630;
        test_addr[993] = 652;
        test_data[993] = 33'd4478315826;
        test_addr[994] = 653;
        test_data[994] = 33'd1452550502;
        test_addr[995] = 654;
        test_data[995] = 33'd3786347631;
        test_addr[996] = 655;
        test_data[996] = 33'd5641215698;
        test_addr[997] = 656;
        test_data[997] = 33'd2873453145;
        test_addr[998] = 657;
        test_data[998] = 33'd5901120262;
        test_addr[999] = 658;
        test_data[999] = 33'd3120144388;
        test_addr[1000] = 659;
        test_data[1000] = 33'd4390205114;
        test_addr[1001] = 660;
        test_data[1001] = 33'd6086763547;
        test_addr[1002] = 661;
        test_data[1002] = 33'd3080712060;
        test_addr[1003] = 527;
        test_data[1003] = 33'd3884199812;
        test_addr[1004] = 528;
        test_data[1004] = 33'd6758356246;
        test_addr[1005] = 529;
        test_data[1005] = 33'd6961602047;
        test_addr[1006] = 530;
        test_data[1006] = 33'd1157531596;
        test_addr[1007] = 531;
        test_data[1007] = 33'd1950799225;
        test_addr[1008] = 532;
        test_data[1008] = 33'd4378687083;
        test_addr[1009] = 533;
        test_data[1009] = 33'd7190073062;
        test_addr[1010] = 771;
        test_data[1010] = 33'd3324619571;
        test_addr[1011] = 772;
        test_data[1011] = 33'd1354814296;
        test_addr[1012] = 773;
        test_data[1012] = 33'd6916470189;
        test_addr[1013] = 774;
        test_data[1013] = 33'd3061105897;
        test_addr[1014] = 775;
        test_data[1014] = 33'd2078638802;
        test_addr[1015] = 776;
        test_data[1015] = 33'd3351180924;
        test_addr[1016] = 777;
        test_data[1016] = 33'd6236484812;
        test_addr[1017] = 778;
        test_data[1017] = 33'd840840300;
        test_addr[1018] = 779;
        test_data[1018] = 33'd1735230795;
        test_addr[1019] = 780;
        test_data[1019] = 33'd7729695326;
        test_addr[1020] = 781;
        test_data[1020] = 33'd7491682468;
        test_addr[1021] = 782;
        test_data[1021] = 33'd4291708288;
        test_addr[1022] = 783;
        test_data[1022] = 33'd655375125;
        test_addr[1023] = 784;
        test_data[1023] = 33'd5058176514;
        test_addr[1024] = 785;
        test_data[1024] = 33'd2189076806;
        test_addr[1025] = 786;
        test_data[1025] = 33'd6141612778;
        test_addr[1026] = 787;
        test_data[1026] = 33'd1740242997;
        test_addr[1027] = 788;
        test_data[1027] = 33'd7687076757;
        test_addr[1028] = 789;
        test_data[1028] = 33'd1888095334;
        test_addr[1029] = 790;
        test_data[1029] = 33'd7975719669;
        test_addr[1030] = 791;
        test_data[1030] = 33'd1151411794;
        test_addr[1031] = 792;
        test_data[1031] = 33'd8187058221;
        test_addr[1032] = 793;
        test_data[1032] = 33'd2283002408;
        test_addr[1033] = 794;
        test_data[1033] = 33'd6507817289;
        test_addr[1034] = 534;
        test_data[1034] = 33'd2544290285;
        test_addr[1035] = 535;
        test_data[1035] = 33'd1551618470;
        test_addr[1036] = 165;
        test_data[1036] = 33'd3597588474;
        test_addr[1037] = 166;
        test_data[1037] = 33'd2253906058;
        test_addr[1038] = 167;
        test_data[1038] = 33'd367704174;
        test_addr[1039] = 168;
        test_data[1039] = 33'd864052885;
        test_addr[1040] = 169;
        test_data[1040] = 33'd7315865421;
        test_addr[1041] = 536;
        test_data[1041] = 33'd6486885970;
        test_addr[1042] = 537;
        test_data[1042] = 33'd1269482248;
        test_addr[1043] = 538;
        test_data[1043] = 33'd2662158238;
        test_addr[1044] = 539;
        test_data[1044] = 33'd1252831804;
        test_addr[1045] = 540;
        test_data[1045] = 33'd3769408227;
        test_addr[1046] = 541;
        test_data[1046] = 33'd6195389909;
        test_addr[1047] = 542;
        test_data[1047] = 33'd5648987651;
        test_addr[1048] = 543;
        test_data[1048] = 33'd108826463;
        test_addr[1049] = 544;
        test_data[1049] = 33'd6794602109;
        test_addr[1050] = 545;
        test_data[1050] = 33'd5988783459;
        test_addr[1051] = 546;
        test_data[1051] = 33'd3953366411;
        test_addr[1052] = 547;
        test_data[1052] = 33'd7078908495;
        test_addr[1053] = 548;
        test_data[1053] = 33'd924290257;
        test_addr[1054] = 549;
        test_data[1054] = 33'd6409850468;
        test_addr[1055] = 550;
        test_data[1055] = 33'd828402464;
        test_addr[1056] = 551;
        test_data[1056] = 33'd3755615061;
        test_addr[1057] = 552;
        test_data[1057] = 33'd2229852656;
        test_addr[1058] = 553;
        test_data[1058] = 33'd3462769718;
        test_addr[1059] = 554;
        test_data[1059] = 33'd5012609015;
        test_addr[1060] = 555;
        test_data[1060] = 33'd3459416445;
        test_addr[1061] = 556;
        test_data[1061] = 33'd2229379164;
        test_addr[1062] = 557;
        test_data[1062] = 33'd6356391616;
        test_addr[1063] = 558;
        test_data[1063] = 33'd1593008829;
        test_addr[1064] = 144;
        test_data[1064] = 33'd1365519167;
        test_addr[1065] = 559;
        test_data[1065] = 33'd1691044550;
        test_addr[1066] = 560;
        test_data[1066] = 33'd2338900121;
        test_addr[1067] = 561;
        test_data[1067] = 33'd5657115115;
        test_addr[1068] = 562;
        test_data[1068] = 33'd3011983409;
        test_addr[1069] = 563;
        test_data[1069] = 33'd3434699751;
        test_addr[1070] = 564;
        test_data[1070] = 33'd869541130;
        test_addr[1071] = 489;
        test_data[1071] = 33'd654573334;
        test_addr[1072] = 490;
        test_data[1072] = 33'd4090258182;
        test_addr[1073] = 491;
        test_data[1073] = 33'd2199790567;
        test_addr[1074] = 492;
        test_data[1074] = 33'd2583156540;
        test_addr[1075] = 493;
        test_data[1075] = 33'd7175925429;
        test_addr[1076] = 494;
        test_data[1076] = 33'd5637581862;
        test_addr[1077] = 495;
        test_data[1077] = 33'd8048378439;
        test_addr[1078] = 496;
        test_data[1078] = 33'd3037540200;
        test_addr[1079] = 497;
        test_data[1079] = 33'd3663618438;
        test_addr[1080] = 498;
        test_data[1080] = 33'd4163492510;
        test_addr[1081] = 499;
        test_data[1081] = 33'd1056200073;
        test_addr[1082] = 500;
        test_data[1082] = 33'd5821379749;
        test_addr[1083] = 501;
        test_data[1083] = 33'd2592532499;
        test_addr[1084] = 502;
        test_data[1084] = 33'd1661402023;
        test_addr[1085] = 565;
        test_data[1085] = 33'd6009749636;
        test_addr[1086] = 566;
        test_data[1086] = 33'd6598486550;
        test_addr[1087] = 567;
        test_data[1087] = 33'd3976280151;
        test_addr[1088] = 568;
        test_data[1088] = 33'd7346398773;
        test_addr[1089] = 569;
        test_data[1089] = 33'd564411764;
        test_addr[1090] = 570;
        test_data[1090] = 33'd4180903970;
        test_addr[1091] = 571;
        test_data[1091] = 33'd3848479732;
        test_addr[1092] = 572;
        test_data[1092] = 33'd403146832;
        test_addr[1093] = 573;
        test_data[1093] = 33'd660266423;
        test_addr[1094] = 574;
        test_data[1094] = 33'd4096603703;
        test_addr[1095] = 575;
        test_data[1095] = 33'd522515645;
        test_addr[1096] = 576;
        test_data[1096] = 33'd8358513562;
        test_addr[1097] = 577;
        test_data[1097] = 33'd469589016;
        test_addr[1098] = 578;
        test_data[1098] = 33'd3176129940;
        test_addr[1099] = 579;
        test_data[1099] = 33'd2815817156;
        test_addr[1100] = 580;
        test_data[1100] = 33'd6981871053;
        test_addr[1101] = 581;
        test_data[1101] = 33'd483805297;
        test_addr[1102] = 582;
        test_data[1102] = 33'd1239020060;
        test_addr[1103] = 583;
        test_data[1103] = 33'd3440524923;
        test_addr[1104] = 584;
        test_data[1104] = 33'd3939647983;
        test_addr[1105] = 585;
        test_data[1105] = 33'd5878626697;
        test_addr[1106] = 586;
        test_data[1106] = 33'd2066734253;
        test_addr[1107] = 587;
        test_data[1107] = 33'd1101126375;
        test_addr[1108] = 588;
        test_data[1108] = 33'd3233337789;
        test_addr[1109] = 589;
        test_data[1109] = 33'd2182645025;
        test_addr[1110] = 590;
        test_data[1110] = 33'd8371970911;
        test_addr[1111] = 591;
        test_data[1111] = 33'd7188573901;
        test_addr[1112] = 592;
        test_data[1112] = 33'd2408379302;
        test_addr[1113] = 593;
        test_data[1113] = 33'd1070801901;
        test_addr[1114] = 594;
        test_data[1114] = 33'd2967625901;
        test_addr[1115] = 595;
        test_data[1115] = 33'd1646515767;
        test_addr[1116] = 596;
        test_data[1116] = 33'd6267662327;
        test_addr[1117] = 597;
        test_data[1117] = 33'd3535940700;
        test_addr[1118] = 598;
        test_data[1118] = 33'd1688883665;
        test_addr[1119] = 328;
        test_data[1119] = 33'd77460711;
        test_addr[1120] = 329;
        test_data[1120] = 33'd6604956318;
        test_addr[1121] = 599;
        test_data[1121] = 33'd6697989393;
        test_addr[1122] = 600;
        test_data[1122] = 33'd4308701688;
        test_addr[1123] = 601;
        test_data[1123] = 33'd1061024359;
        test_addr[1124] = 602;
        test_data[1124] = 33'd7935273800;
        test_addr[1125] = 603;
        test_data[1125] = 33'd7087584803;
        test_addr[1126] = 604;
        test_data[1126] = 33'd1113088347;
        test_addr[1127] = 605;
        test_data[1127] = 33'd1618144234;
        test_addr[1128] = 606;
        test_data[1128] = 33'd920782161;
        test_addr[1129] = 390;
        test_data[1129] = 33'd2543760664;
        test_addr[1130] = 391;
        test_data[1130] = 33'd189757725;
        test_addr[1131] = 392;
        test_data[1131] = 33'd1006684681;
        test_addr[1132] = 393;
        test_data[1132] = 33'd479449245;
        test_addr[1133] = 394;
        test_data[1133] = 33'd7726484703;
        test_addr[1134] = 395;
        test_data[1134] = 33'd6030052594;
        test_addr[1135] = 396;
        test_data[1135] = 33'd5195098441;
        test_addr[1136] = 397;
        test_data[1136] = 33'd4140998441;
        test_addr[1137] = 398;
        test_data[1137] = 33'd3505084960;
        test_addr[1138] = 399;
        test_data[1138] = 33'd1244846146;
        test_addr[1139] = 400;
        test_data[1139] = 33'd5806859320;
        test_addr[1140] = 607;
        test_data[1140] = 33'd3986635328;
        test_addr[1141] = 608;
        test_data[1141] = 33'd2953791377;
        test_addr[1142] = 609;
        test_data[1142] = 33'd3511563354;
        test_addr[1143] = 610;
        test_data[1143] = 33'd2559326217;
        test_addr[1144] = 611;
        test_data[1144] = 33'd2941323753;
        test_addr[1145] = 612;
        test_data[1145] = 33'd8001268366;
        test_addr[1146] = 613;
        test_data[1146] = 33'd5365713684;
        test_addr[1147] = 614;
        test_data[1147] = 33'd2106134210;
        test_addr[1148] = 615;
        test_data[1148] = 33'd4288664088;
        test_addr[1149] = 616;
        test_data[1149] = 33'd6574817601;
        test_addr[1150] = 617;
        test_data[1150] = 33'd1884511967;
        test_addr[1151] = 618;
        test_data[1151] = 33'd7004053359;
        test_addr[1152] = 619;
        test_data[1152] = 33'd7434932244;
        test_addr[1153] = 620;
        test_data[1153] = 33'd2147528937;
        test_addr[1154] = 621;
        test_data[1154] = 33'd765391404;
        test_addr[1155] = 622;
        test_data[1155] = 33'd6784844864;
        test_addr[1156] = 623;
        test_data[1156] = 33'd2373385250;
        test_addr[1157] = 624;
        test_data[1157] = 33'd8315716912;
        test_addr[1158] = 625;
        test_data[1158] = 33'd1909344899;
        test_addr[1159] = 626;
        test_data[1159] = 33'd3411209394;
        test_addr[1160] = 627;
        test_data[1160] = 33'd111369000;
        test_addr[1161] = 628;
        test_data[1161] = 33'd108823116;
        test_addr[1162] = 629;
        test_data[1162] = 33'd4225840529;
        test_addr[1163] = 630;
        test_data[1163] = 33'd911457724;
        test_addr[1164] = 631;
        test_data[1164] = 33'd4116914749;
        test_addr[1165] = 632;
        test_data[1165] = 33'd5588247199;
        test_addr[1166] = 633;
        test_data[1166] = 33'd1090431518;
        test_addr[1167] = 966;
        test_data[1167] = 33'd2186720106;
        test_addr[1168] = 967;
        test_data[1168] = 33'd227677533;
        test_addr[1169] = 968;
        test_data[1169] = 33'd6979391612;
        test_addr[1170] = 969;
        test_data[1170] = 33'd7874843620;
        test_addr[1171] = 970;
        test_data[1171] = 33'd2846411311;
        test_addr[1172] = 971;
        test_data[1172] = 33'd7316913241;
        test_addr[1173] = 972;
        test_data[1173] = 33'd3134925533;
        test_addr[1174] = 973;
        test_data[1174] = 33'd2724948106;
        test_addr[1175] = 974;
        test_data[1175] = 33'd6858535231;
        test_addr[1176] = 975;
        test_data[1176] = 33'd267738865;
        test_addr[1177] = 634;
        test_data[1177] = 33'd3651902078;
        test_addr[1178] = 455;
        test_data[1178] = 33'd6642941137;
        test_addr[1179] = 456;
        test_data[1179] = 33'd2010861474;
        test_addr[1180] = 457;
        test_data[1180] = 33'd15769730;
        test_addr[1181] = 635;
        test_data[1181] = 33'd3605989952;
        test_addr[1182] = 636;
        test_data[1182] = 33'd1964111665;
        test_addr[1183] = 637;
        test_data[1183] = 33'd4716483905;
        test_addr[1184] = 638;
        test_data[1184] = 33'd3568991821;
        test_addr[1185] = 639;
        test_data[1185] = 33'd4062177817;
        test_addr[1186] = 640;
        test_data[1186] = 33'd3889086438;
        test_addr[1187] = 641;
        test_data[1187] = 33'd3812820741;
        test_addr[1188] = 233;
        test_data[1188] = 33'd2492348860;
        test_addr[1189] = 234;
        test_data[1189] = 33'd3059098805;
        test_addr[1190] = 235;
        test_data[1190] = 33'd379016448;
        test_addr[1191] = 236;
        test_data[1191] = 33'd6548423851;
        test_addr[1192] = 237;
        test_data[1192] = 33'd3293190254;
        test_addr[1193] = 238;
        test_data[1193] = 33'd7018267365;
        test_addr[1194] = 239;
        test_data[1194] = 33'd1677771600;
        test_addr[1195] = 240;
        test_data[1195] = 33'd4627671479;
        test_addr[1196] = 241;
        test_data[1196] = 33'd3112036660;
        test_addr[1197] = 242;
        test_data[1197] = 33'd502196391;
        test_addr[1198] = 243;
        test_data[1198] = 33'd1440318250;
        test_addr[1199] = 244;
        test_data[1199] = 33'd1318439210;
        test_addr[1200] = 245;
        test_data[1200] = 33'd324506329;
        test_addr[1201] = 246;
        test_data[1201] = 33'd801919684;
        test_addr[1202] = 247;
        test_data[1202] = 33'd3793934249;
        test_addr[1203] = 642;
        test_data[1203] = 33'd982240008;
        test_addr[1204] = 643;
        test_data[1204] = 33'd5332629428;
        test_addr[1205] = 644;
        test_data[1205] = 33'd3029388123;
        test_addr[1206] = 645;
        test_data[1206] = 33'd199889460;
        test_addr[1207] = 646;
        test_data[1207] = 33'd1325289533;
        test_addr[1208] = 647;
        test_data[1208] = 33'd1303442273;
        test_addr[1209] = 648;
        test_data[1209] = 33'd2300180881;
        test_addr[1210] = 649;
        test_data[1210] = 33'd8480746332;
        test_addr[1211] = 252;
        test_data[1211] = 33'd855026393;
        test_addr[1212] = 253;
        test_data[1212] = 33'd7139286089;
        test_addr[1213] = 254;
        test_data[1213] = 33'd100893370;
        test_addr[1214] = 255;
        test_data[1214] = 33'd3493356248;
        test_addr[1215] = 650;
        test_data[1215] = 33'd7305742169;
        test_addr[1216] = 651;
        test_data[1216] = 33'd7710424776;
        test_addr[1217] = 270;
        test_data[1217] = 33'd4155868294;
        test_addr[1218] = 271;
        test_data[1218] = 33'd1009868606;
        test_addr[1219] = 652;
        test_data[1219] = 33'd183348530;
        test_addr[1220] = 653;
        test_data[1220] = 33'd1452550502;
        test_addr[1221] = 654;
        test_data[1221] = 33'd3786347631;
        test_addr[1222] = 655;
        test_data[1222] = 33'd1346248402;
        test_addr[1223] = 656;
        test_data[1223] = 33'd6870542609;
        test_addr[1224] = 657;
        test_data[1224] = 33'd1606152966;
        test_addr[1225] = 658;
        test_data[1225] = 33'd3120144388;
        test_addr[1226] = 659;
        test_data[1226] = 33'd7480471368;
        test_addr[1227] = 660;
        test_data[1227] = 33'd1791796251;
        test_addr[1228] = 661;
        test_data[1228] = 33'd3080712060;
        test_addr[1229] = 662;
        test_data[1229] = 33'd4978667645;
        test_addr[1230] = 663;
        test_data[1230] = 33'd89312420;
        test_addr[1231] = 664;
        test_data[1231] = 33'd4123313617;
        test_addr[1232] = 665;
        test_data[1232] = 33'd5529169153;
        test_addr[1233] = 666;
        test_data[1233] = 33'd812647693;
        test_addr[1234] = 667;
        test_data[1234] = 33'd560999711;
        test_addr[1235] = 668;
        test_data[1235] = 33'd4073128129;
        test_addr[1236] = 83;
        test_data[1236] = 33'd6827783459;
        test_addr[1237] = 84;
        test_data[1237] = 33'd655204540;
        test_addr[1238] = 85;
        test_data[1238] = 33'd4108519334;
        test_addr[1239] = 86;
        test_data[1239] = 33'd4331752554;
        test_addr[1240] = 87;
        test_data[1240] = 33'd1074381877;
        test_addr[1241] = 88;
        test_data[1241] = 33'd4145639023;
        test_addr[1242] = 89;
        test_data[1242] = 33'd3402301464;
        test_addr[1243] = 90;
        test_data[1243] = 33'd8103868626;
        test_addr[1244] = 91;
        test_data[1244] = 33'd2419969866;
        test_addr[1245] = 92;
        test_data[1245] = 33'd1952513095;
        test_addr[1246] = 93;
        test_data[1246] = 33'd1228061459;
        test_addr[1247] = 669;
        test_data[1247] = 33'd716422625;
        test_addr[1248] = 665;
        test_data[1248] = 33'd1234201857;
        test_addr[1249] = 670;
        test_data[1249] = 33'd8571485769;
        test_addr[1250] = 671;
        test_data[1250] = 33'd2151985146;
        test_addr[1251] = 672;
        test_data[1251] = 33'd7133827392;
        test_addr[1252] = 673;
        test_data[1252] = 33'd2206060871;
        test_addr[1253] = 674;
        test_data[1253] = 33'd5906943610;
        test_addr[1254] = 675;
        test_data[1254] = 33'd3430516374;
        test_addr[1255] = 676;
        test_data[1255] = 33'd662578081;
        test_addr[1256] = 677;
        test_data[1256] = 33'd2331235146;
        test_addr[1257] = 678;
        test_data[1257] = 33'd8497918065;
        test_addr[1258] = 679;
        test_data[1258] = 33'd6602221863;
        test_addr[1259] = 680;
        test_data[1259] = 33'd772379733;
        test_addr[1260] = 681;
        test_data[1260] = 33'd85007220;
        test_addr[1261] = 682;
        test_data[1261] = 33'd666405120;
        test_addr[1262] = 683;
        test_data[1262] = 33'd1731237928;
        test_addr[1263] = 684;
        test_data[1263] = 33'd6476778885;
        test_addr[1264] = 685;
        test_data[1264] = 33'd4976250764;
        test_addr[1265] = 686;
        test_data[1265] = 33'd4109187007;
        test_addr[1266] = 687;
        test_data[1266] = 33'd8099228872;
        test_addr[1267] = 87;
        test_data[1267] = 33'd1074381877;
        test_addr[1268] = 88;
        test_data[1268] = 33'd5857239192;
        test_addr[1269] = 89;
        test_data[1269] = 33'd7561158962;
        test_addr[1270] = 90;
        test_data[1270] = 33'd5142752616;
        test_addr[1271] = 91;
        test_data[1271] = 33'd5145239925;
        test_addr[1272] = 92;
        test_data[1272] = 33'd1952513095;
        test_addr[1273] = 93;
        test_data[1273] = 33'd6519945864;
        test_addr[1274] = 94;
        test_data[1274] = 33'd3836173812;
        test_addr[1275] = 95;
        test_data[1275] = 33'd310852482;
        test_addr[1276] = 96;
        test_data[1276] = 33'd6016149844;
        test_addr[1277] = 97;
        test_data[1277] = 33'd3946323928;
        test_addr[1278] = 98;
        test_data[1278] = 33'd7809852884;
        test_addr[1279] = 99;
        test_data[1279] = 33'd3402368761;
        test_addr[1280] = 100;
        test_data[1280] = 33'd2034825318;
        test_addr[1281] = 101;
        test_data[1281] = 33'd6370518697;
        test_addr[1282] = 102;
        test_data[1282] = 33'd457023927;
        test_addr[1283] = 688;
        test_data[1283] = 33'd2293783707;
        test_addr[1284] = 689;
        test_data[1284] = 33'd2765668052;
        test_addr[1285] = 690;
        test_data[1285] = 33'd4391808570;
        test_addr[1286] = 691;
        test_data[1286] = 33'd7584460848;
        test_addr[1287] = 692;
        test_data[1287] = 33'd984956215;
        test_addr[1288] = 693;
        test_data[1288] = 33'd6371002124;
        test_addr[1289] = 694;
        test_data[1289] = 33'd7631453384;
        test_addr[1290] = 597;
        test_data[1290] = 33'd3535940700;
        test_addr[1291] = 598;
        test_data[1291] = 33'd8406491916;
        test_addr[1292] = 599;
        test_data[1292] = 33'd2403022097;
        test_addr[1293] = 600;
        test_data[1293] = 33'd7379486238;
        test_addr[1294] = 695;
        test_data[1294] = 33'd4659718123;
        test_addr[1295] = 696;
        test_data[1295] = 33'd2824012066;
        test_addr[1296] = 697;
        test_data[1296] = 33'd2908751719;
        test_addr[1297] = 698;
        test_data[1297] = 33'd2093503010;
        test_addr[1298] = 699;
        test_data[1298] = 33'd3070843493;
        test_addr[1299] = 700;
        test_data[1299] = 33'd1020382117;
        test_addr[1300] = 701;
        test_data[1300] = 33'd6184088391;
        test_addr[1301] = 702;
        test_data[1301] = 33'd5432885875;
        test_addr[1302] = 703;
        test_data[1302] = 33'd2023405860;
        test_addr[1303] = 704;
        test_data[1303] = 33'd5471894294;
        test_addr[1304] = 705;
        test_data[1304] = 33'd4570153214;
        test_addr[1305] = 706;
        test_data[1305] = 33'd3602815316;
        test_addr[1306] = 707;
        test_data[1306] = 33'd3409958362;
        test_addr[1307] = 708;
        test_data[1307] = 33'd3004227477;
        test_addr[1308] = 709;
        test_data[1308] = 33'd265858089;
        test_addr[1309] = 710;
        test_data[1309] = 33'd868282533;
        test_addr[1310] = 711;
        test_data[1310] = 33'd8019391752;
        test_addr[1311] = 567;
        test_data[1311] = 33'd3976280151;
        test_addr[1312] = 568;
        test_data[1312] = 33'd5731039904;
        test_addr[1313] = 569;
        test_data[1313] = 33'd5819918080;
        test_addr[1314] = 712;
        test_data[1314] = 33'd6755060679;
        test_addr[1315] = 713;
        test_data[1315] = 33'd4466036316;
        test_addr[1316] = 714;
        test_data[1316] = 33'd299549045;
        test_addr[1317] = 715;
        test_data[1317] = 33'd6820531657;
        test_addr[1318] = 716;
        test_data[1318] = 33'd292650974;
        test_addr[1319] = 717;
        test_data[1319] = 33'd5565228692;
        test_addr[1320] = 718;
        test_data[1320] = 33'd3656605274;
        test_addr[1321] = 719;
        test_data[1321] = 33'd5608232235;
        test_addr[1322] = 720;
        test_data[1322] = 33'd264781874;
        test_addr[1323] = 721;
        test_data[1323] = 33'd579303093;
        test_addr[1324] = 722;
        test_data[1324] = 33'd1583494039;
        test_addr[1325] = 723;
        test_data[1325] = 33'd7855165078;
        test_addr[1326] = 724;
        test_data[1326] = 33'd1061855659;
        test_addr[1327] = 725;
        test_data[1327] = 33'd7581709874;
        test_addr[1328] = 726;
        test_data[1328] = 33'd8512437101;
        test_addr[1329] = 727;
        test_data[1329] = 33'd2678040300;
        test_addr[1330] = 728;
        test_data[1330] = 33'd2822296548;
        test_addr[1331] = 729;
        test_data[1331] = 33'd578785750;
        test_addr[1332] = 227;
        test_data[1332] = 33'd2688484918;
        test_addr[1333] = 228;
        test_data[1333] = 33'd4120475529;
        test_addr[1334] = 229;
        test_data[1334] = 33'd665005425;
        test_addr[1335] = 230;
        test_data[1335] = 33'd988458485;
        test_addr[1336] = 231;
        test_data[1336] = 33'd2346487764;
        test_addr[1337] = 232;
        test_data[1337] = 33'd5959996415;
        test_addr[1338] = 233;
        test_data[1338] = 33'd2492348860;
        test_addr[1339] = 234;
        test_data[1339] = 33'd3059098805;
        test_addr[1340] = 235;
        test_data[1340] = 33'd4892522500;
        test_addr[1341] = 236;
        test_data[1341] = 33'd2253456555;
        test_addr[1342] = 237;
        test_data[1342] = 33'd5149264602;
        test_addr[1343] = 238;
        test_data[1343] = 33'd2723300069;
        test_addr[1344] = 239;
        test_data[1344] = 33'd1677771600;
        test_addr[1345] = 730;
        test_data[1345] = 33'd2998442618;
        test_addr[1346] = 731;
        test_data[1346] = 33'd6579830709;
        test_addr[1347] = 732;
        test_data[1347] = 33'd1766000469;
        test_addr[1348] = 733;
        test_data[1348] = 33'd3548136803;
        test_addr[1349] = 734;
        test_data[1349] = 33'd1311988770;
        test_addr[1350] = 735;
        test_data[1350] = 33'd3996876697;
        test_addr[1351] = 242;
        test_data[1351] = 33'd502196391;
        test_addr[1352] = 243;
        test_data[1352] = 33'd7778424111;
        test_addr[1353] = 244;
        test_data[1353] = 33'd1318439210;
        test_addr[1354] = 245;
        test_data[1354] = 33'd324506329;
        test_addr[1355] = 736;
        test_data[1355] = 33'd3833161201;
        test_addr[1356] = 737;
        test_data[1356] = 33'd4894420229;
        test_addr[1357] = 738;
        test_data[1357] = 33'd5857784515;
        test_addr[1358] = 739;
        test_data[1358] = 33'd6876160315;
        test_addr[1359] = 740;
        test_data[1359] = 33'd725439312;
        test_addr[1360] = 741;
        test_data[1360] = 33'd336889000;
        test_addr[1361] = 742;
        test_data[1361] = 33'd5985466922;
        test_addr[1362] = 743;
        test_data[1362] = 33'd3044130341;
        test_addr[1363] = 744;
        test_data[1363] = 33'd1292464610;
        test_addr[1364] = 745;
        test_data[1364] = 33'd4084688614;
        test_addr[1365] = 746;
        test_data[1365] = 33'd689947192;
        test_addr[1366] = 747;
        test_data[1366] = 33'd4343687905;
        test_addr[1367] = 748;
        test_data[1367] = 33'd76408912;
        test_addr[1368] = 749;
        test_data[1368] = 33'd821619415;
        test_addr[1369] = 750;
        test_data[1369] = 33'd1056728340;
        test_addr[1370] = 751;
        test_data[1370] = 33'd6950207487;
        test_addr[1371] = 752;
        test_data[1371] = 33'd8048822140;
        test_addr[1372] = 753;
        test_data[1372] = 33'd5589627859;
        test_addr[1373] = 754;
        test_data[1373] = 33'd1731907904;
        test_addr[1374] = 755;
        test_data[1374] = 33'd1320792984;
        test_addr[1375] = 756;
        test_data[1375] = 33'd2829182134;
        test_addr[1376] = 757;
        test_data[1376] = 33'd5523480713;
        test_addr[1377] = 758;
        test_data[1377] = 33'd3678702924;
        test_addr[1378] = 759;
        test_data[1378] = 33'd3506733921;
        test_addr[1379] = 760;
        test_data[1379] = 33'd3222496793;
        test_addr[1380] = 761;
        test_data[1380] = 33'd813817359;
        test_addr[1381] = 762;
        test_data[1381] = 33'd8523184784;
        test_addr[1382] = 763;
        test_data[1382] = 33'd407903955;
        test_addr[1383] = 764;
        test_data[1383] = 33'd5139013858;
        test_addr[1384] = 765;
        test_data[1384] = 33'd8410563357;
        test_addr[1385] = 766;
        test_data[1385] = 33'd7241747587;
        test_addr[1386] = 48;
        test_data[1386] = 33'd4413986114;
        test_addr[1387] = 49;
        test_data[1387] = 33'd3795521150;
        test_addr[1388] = 50;
        test_data[1388] = 33'd4466023831;
        test_addr[1389] = 51;
        test_data[1389] = 33'd3965955358;
        test_addr[1390] = 52;
        test_data[1390] = 33'd1670309798;
        test_addr[1391] = 53;
        test_data[1391] = 33'd5665899954;
        test_addr[1392] = 54;
        test_data[1392] = 33'd3762196439;
        test_addr[1393] = 55;
        test_data[1393] = 33'd3541808763;
        test_addr[1394] = 56;
        test_data[1394] = 33'd4032767092;
        test_addr[1395] = 57;
        test_data[1395] = 33'd3015078990;
        test_addr[1396] = 58;
        test_data[1396] = 33'd2630100688;
        test_addr[1397] = 767;
        test_data[1397] = 33'd51594790;
        test_addr[1398] = 768;
        test_data[1398] = 33'd2995316459;
        test_addr[1399] = 769;
        test_data[1399] = 33'd2466504171;
        test_addr[1400] = 770;
        test_data[1400] = 33'd8470092981;
        test_addr[1401] = 771;
        test_data[1401] = 33'd3324619571;
        test_addr[1402] = 772;
        test_data[1402] = 33'd1354814296;
        test_addr[1403] = 773;
        test_data[1403] = 33'd2621502893;
        test_addr[1404] = 774;
        test_data[1404] = 33'd3061105897;
        test_addr[1405] = 775;
        test_data[1405] = 33'd7261749658;
        test_addr[1406] = 854;
        test_data[1406] = 33'd2265029546;
        test_addr[1407] = 855;
        test_data[1407] = 33'd325563839;
        test_addr[1408] = 856;
        test_data[1408] = 33'd1518218722;
        test_addr[1409] = 857;
        test_data[1409] = 33'd456204038;
        test_addr[1410] = 858;
        test_data[1410] = 33'd2316112060;
        test_addr[1411] = 859;
        test_data[1411] = 33'd8291181225;
        test_addr[1412] = 860;
        test_data[1412] = 33'd9740189;
        test_addr[1413] = 861;
        test_data[1413] = 33'd6906712573;
        test_addr[1414] = 862;
        test_data[1414] = 33'd6186141872;
        test_addr[1415] = 863;
        test_data[1415] = 33'd3181973309;
        test_addr[1416] = 864;
        test_data[1416] = 33'd5970539606;
        test_addr[1417] = 865;
        test_data[1417] = 33'd2442557656;
        test_addr[1418] = 866;
        test_data[1418] = 33'd6920341800;
        test_addr[1419] = 867;
        test_data[1419] = 33'd4191967086;
        test_addr[1420] = 868;
        test_data[1420] = 33'd7914255644;
        test_addr[1421] = 869;
        test_data[1421] = 33'd7570366732;
        test_addr[1422] = 870;
        test_data[1422] = 33'd747559002;
        test_addr[1423] = 871;
        test_data[1423] = 33'd5395256937;
        test_addr[1424] = 872;
        test_data[1424] = 33'd3833194746;
        test_addr[1425] = 873;
        test_data[1425] = 33'd1130221406;
        test_addr[1426] = 776;
        test_data[1426] = 33'd3351180924;
        test_addr[1427] = 777;
        test_data[1427] = 33'd1941517516;
        test_addr[1428] = 778;
        test_data[1428] = 33'd7953471692;
        test_addr[1429] = 120;
        test_data[1429] = 33'd2264552573;
        test_addr[1430] = 121;
        test_data[1430] = 33'd2605200182;
        test_addr[1431] = 122;
        test_data[1431] = 33'd3622924683;
        test_addr[1432] = 123;
        test_data[1432] = 33'd5754524903;
        test_addr[1433] = 124;
        test_data[1433] = 33'd386667355;
        test_addr[1434] = 125;
        test_data[1434] = 33'd1182003256;
        test_addr[1435] = 126;
        test_data[1435] = 33'd989367641;
        test_addr[1436] = 127;
        test_data[1436] = 33'd5267767702;
        test_addr[1437] = 128;
        test_data[1437] = 33'd2116858368;
        test_addr[1438] = 129;
        test_data[1438] = 33'd212359631;
        test_addr[1439] = 130;
        test_data[1439] = 33'd3185392084;
        test_addr[1440] = 131;
        test_data[1440] = 33'd2412978687;
        test_addr[1441] = 779;
        test_data[1441] = 33'd1735230795;
        test_addr[1442] = 780;
        test_data[1442] = 33'd3434728030;
        test_addr[1443] = 781;
        test_data[1443] = 33'd7027657595;
        test_addr[1444] = 782;
        test_data[1444] = 33'd4291708288;
        test_addr[1445] = 783;
        test_data[1445] = 33'd655375125;
        test_addr[1446] = 784;
        test_data[1446] = 33'd5889748662;
        test_addr[1447] = 785;
        test_data[1447] = 33'd2189076806;
        test_addr[1448] = 786;
        test_data[1448] = 33'd5069974466;
        test_addr[1449] = 787;
        test_data[1449] = 33'd1740242997;
        test_addr[1450] = 788;
        test_data[1450] = 33'd3392109461;
        test_addr[1451] = 789;
        test_data[1451] = 33'd1888095334;
        test_addr[1452] = 790;
        test_data[1452] = 33'd3680752373;
        test_addr[1453] = 791;
        test_data[1453] = 33'd1151411794;
        test_addr[1454] = 792;
        test_data[1454] = 33'd7585232240;
        test_addr[1455] = 793;
        test_data[1455] = 33'd2283002408;
        test_addr[1456] = 843;
        test_data[1456] = 33'd3444648562;
        test_addr[1457] = 844;
        test_data[1457] = 33'd7921379097;
        test_addr[1458] = 845;
        test_data[1458] = 33'd7043772286;
        test_addr[1459] = 846;
        test_data[1459] = 33'd3129315442;
        test_addr[1460] = 847;
        test_data[1460] = 33'd1929108195;
        test_addr[1461] = 848;
        test_data[1461] = 33'd2055262394;
        test_addr[1462] = 849;
        test_data[1462] = 33'd8555245157;
        test_addr[1463] = 850;
        test_data[1463] = 33'd1598966603;
        test_addr[1464] = 851;
        test_data[1464] = 33'd5343335175;
        test_addr[1465] = 794;
        test_data[1465] = 33'd2212849993;
        test_addr[1466] = 795;
        test_data[1466] = 33'd2128607902;
        test_addr[1467] = 796;
        test_data[1467] = 33'd4275211649;
        test_addr[1468] = 797;
        test_data[1468] = 33'd3562187736;
        test_addr[1469] = 798;
        test_data[1469] = 33'd4098353399;
        test_addr[1470] = 799;
        test_data[1470] = 33'd1518077955;
        test_addr[1471] = 800;
        test_data[1471] = 33'd754500382;
        test_addr[1472] = 801;
        test_data[1472] = 33'd584393855;
        test_addr[1473] = 802;
        test_data[1473] = 33'd3063225216;
        test_addr[1474] = 803;
        test_data[1474] = 33'd1034772483;
        test_addr[1475] = 804;
        test_data[1475] = 33'd8294198066;
        test_addr[1476] = 805;
        test_data[1476] = 33'd2518139456;
        test_addr[1477] = 806;
        test_data[1477] = 33'd1466474561;
        test_addr[1478] = 807;
        test_data[1478] = 33'd639577463;
        test_addr[1479] = 316;
        test_data[1479] = 33'd498221104;
        test_addr[1480] = 317;
        test_data[1480] = 33'd2374556068;
        test_addr[1481] = 318;
        test_data[1481] = 33'd2835077050;
        test_addr[1482] = 319;
        test_data[1482] = 33'd357113237;
        test_addr[1483] = 320;
        test_data[1483] = 33'd2364460379;
        test_addr[1484] = 321;
        test_data[1484] = 33'd8573947021;
        test_addr[1485] = 322;
        test_data[1485] = 33'd341336502;
        test_addr[1486] = 323;
        test_data[1486] = 33'd6248766529;
        test_addr[1487] = 324;
        test_data[1487] = 33'd6409771942;
        test_addr[1488] = 325;
        test_data[1488] = 33'd2617615466;
        test_addr[1489] = 326;
        test_data[1489] = 33'd4881430980;
        test_addr[1490] = 327;
        test_data[1490] = 33'd739327056;
        test_addr[1491] = 328;
        test_data[1491] = 33'd7203333425;
        test_addr[1492] = 329;
        test_data[1492] = 33'd2309989022;
        test_addr[1493] = 330;
        test_data[1493] = 33'd3508612389;
        test_addr[1494] = 331;
        test_data[1494] = 33'd4229591735;
        test_addr[1495] = 332;
        test_data[1495] = 33'd4266769130;
        test_addr[1496] = 808;
        test_data[1496] = 33'd8459002353;
        test_addr[1497] = 809;
        test_data[1497] = 33'd3968329823;
        test_addr[1498] = 810;
        test_data[1498] = 33'd5963120298;
        test_addr[1499] = 811;
        test_data[1499] = 33'd2968812544;
        test_addr[1500] = 812;
        test_data[1500] = 33'd7239596612;
        test_addr[1501] = 813;
        test_data[1501] = 33'd3207399348;
        test_addr[1502] = 566;
        test_data[1502] = 33'd2303519254;
        test_addr[1503] = 567;
        test_data[1503] = 33'd3976280151;
        test_addr[1504] = 568;
        test_data[1504] = 33'd7662060043;
        test_addr[1505] = 569;
        test_data[1505] = 33'd1524950784;
        test_addr[1506] = 570;
        test_data[1506] = 33'd4180903970;
        test_addr[1507] = 571;
        test_data[1507] = 33'd3848479732;
        test_addr[1508] = 572;
        test_data[1508] = 33'd403146832;
        test_addr[1509] = 573;
        test_data[1509] = 33'd660266423;
        test_addr[1510] = 574;
        test_data[1510] = 33'd7490582948;
        test_addr[1511] = 575;
        test_data[1511] = 33'd522515645;
        test_addr[1512] = 576;
        test_data[1512] = 33'd4644735780;
        test_addr[1513] = 577;
        test_data[1513] = 33'd469589016;
        test_addr[1514] = 578;
        test_data[1514] = 33'd3176129940;
        test_addr[1515] = 579;
        test_data[1515] = 33'd2815817156;
        test_addr[1516] = 580;
        test_data[1516] = 33'd2686903757;
        test_addr[1517] = 581;
        test_data[1517] = 33'd483805297;
        test_addr[1518] = 814;
        test_data[1518] = 33'd2532614522;
        test_addr[1519] = 815;
        test_data[1519] = 33'd7891433285;
        test_addr[1520] = 816;
        test_data[1520] = 33'd2089907260;
        test_addr[1521] = 817;
        test_data[1521] = 33'd7834135682;
        test_addr[1522] = 818;
        test_data[1522] = 33'd7430106334;
        test_addr[1523] = 819;
        test_data[1523] = 33'd3407332409;
        test_addr[1524] = 820;
        test_data[1524] = 33'd3200758228;
        test_addr[1525] = 821;
        test_data[1525] = 33'd131890680;
        test_addr[1526] = 822;
        test_data[1526] = 33'd2790105153;
        test_addr[1527] = 823;
        test_data[1527] = 33'd6236560545;
        test_addr[1528] = 824;
        test_data[1528] = 33'd4185437212;
        test_addr[1529] = 825;
        test_data[1529] = 33'd1444494147;
        test_addr[1530] = 826;
        test_data[1530] = 33'd4588799873;
        test_addr[1531] = 827;
        test_data[1531] = 33'd4271161680;
        test_addr[1532] = 828;
        test_data[1532] = 33'd8523434429;
        test_addr[1533] = 580;
        test_data[1533] = 33'd2686903757;
        test_addr[1534] = 581;
        test_data[1534] = 33'd483805297;
        test_addr[1535] = 582;
        test_data[1535] = 33'd4856297806;
        test_addr[1536] = 829;
        test_data[1536] = 33'd2471067861;
        test_addr[1537] = 830;
        test_data[1537] = 33'd2151514164;
        test_addr[1538] = 831;
        test_data[1538] = 33'd3512387836;
        test_addr[1539] = 832;
        test_data[1539] = 33'd2442866266;
        test_addr[1540] = 833;
        test_data[1540] = 33'd6052184422;
        test_addr[1541] = 880;
        test_data[1541] = 33'd1009940429;
        test_addr[1542] = 834;
        test_data[1542] = 33'd1624961981;
        test_addr[1543] = 835;
        test_data[1543] = 33'd3185900460;
        test_addr[1544] = 836;
        test_data[1544] = 33'd2868439311;
        test_addr[1545] = 837;
        test_data[1545] = 33'd6589978914;
        test_addr[1546] = 838;
        test_data[1546] = 33'd2598268969;
        test_addr[1547] = 839;
        test_data[1547] = 33'd2544945082;
        test_addr[1548] = 840;
        test_data[1548] = 33'd2690967453;
        test_addr[1549] = 841;
        test_data[1549] = 33'd3495259579;
        test_addr[1550] = 842;
        test_data[1550] = 33'd6216360960;
        test_addr[1551] = 843;
        test_data[1551] = 33'd3444648562;
        test_addr[1552] = 844;
        test_data[1552] = 33'd5199445551;
        test_addr[1553] = 845;
        test_data[1553] = 33'd2748804990;
        test_addr[1554] = 846;
        test_data[1554] = 33'd3129315442;
        test_addr[1555] = 847;
        test_data[1555] = 33'd1929108195;
        test_addr[1556] = 848;
        test_data[1556] = 33'd2055262394;
        test_addr[1557] = 849;
        test_data[1557] = 33'd4260277861;
        test_addr[1558] = 850;
        test_data[1558] = 33'd1598966603;
        test_addr[1559] = 851;
        test_data[1559] = 33'd1048367879;
        test_addr[1560] = 852;
        test_data[1560] = 33'd4396436069;
        test_addr[1561] = 853;
        test_data[1561] = 33'd1560350512;
        test_addr[1562] = 854;
        test_data[1562] = 33'd7626911191;
        test_addr[1563] = 855;
        test_data[1563] = 33'd5562579323;
        test_addr[1564] = 856;
        test_data[1564] = 33'd6291504930;
        test_addr[1565] = 857;
        test_data[1565] = 33'd5345753294;
        test_addr[1566] = 858;
        test_data[1566] = 33'd5892266000;
        test_addr[1567] = 859;
        test_data[1567] = 33'd3996213929;
        test_addr[1568] = 860;
        test_data[1568] = 33'd9740189;
        test_addr[1569] = 861;
        test_data[1569] = 33'd2611745277;
        test_addr[1570] = 428;
        test_data[1570] = 33'd807619004;
        test_addr[1571] = 429;
        test_data[1571] = 33'd4094634244;
        test_addr[1572] = 430;
        test_data[1572] = 33'd896214945;
        test_addr[1573] = 431;
        test_data[1573] = 33'd3279784998;
        test_addr[1574] = 432;
        test_data[1574] = 33'd842198295;
        test_addr[1575] = 433;
        test_data[1575] = 33'd1529853911;
        test_addr[1576] = 434;
        test_data[1576] = 33'd423001153;
        test_addr[1577] = 435;
        test_data[1577] = 33'd2315575124;
        test_addr[1578] = 436;
        test_data[1578] = 33'd4034103201;
        test_addr[1579] = 437;
        test_data[1579] = 33'd2303126498;
        test_addr[1580] = 438;
        test_data[1580] = 33'd6150919642;
        test_addr[1581] = 439;
        test_data[1581] = 33'd3187307611;
        test_addr[1582] = 440;
        test_data[1582] = 33'd731387276;
        test_addr[1583] = 441;
        test_data[1583] = 33'd2079610815;
        test_addr[1584] = 442;
        test_data[1584] = 33'd4928209920;
        test_addr[1585] = 443;
        test_data[1585] = 33'd8498956342;
        test_addr[1586] = 444;
        test_data[1586] = 33'd2677223067;
        test_addr[1587] = 445;
        test_data[1587] = 33'd637046458;
        test_addr[1588] = 446;
        test_data[1588] = 33'd1320511667;
        test_addr[1589] = 447;
        test_data[1589] = 33'd3084548448;
        test_addr[1590] = 448;
        test_data[1590] = 33'd2047532963;
        test_addr[1591] = 449;
        test_data[1591] = 33'd658651725;
        test_addr[1592] = 450;
        test_data[1592] = 33'd8584870185;
        test_addr[1593] = 451;
        test_data[1593] = 33'd772375377;
        test_addr[1594] = 452;
        test_data[1594] = 33'd1012981055;
        test_addr[1595] = 453;
        test_data[1595] = 33'd4144249236;
        test_addr[1596] = 454;
        test_data[1596] = 33'd3006483553;
        test_addr[1597] = 455;
        test_data[1597] = 33'd7775869411;
        test_addr[1598] = 456;
        test_data[1598] = 33'd2010861474;
        test_addr[1599] = 457;
        test_data[1599] = 33'd15769730;
        test_addr[1600] = 862;
        test_data[1600] = 33'd5664522208;
        test_addr[1601] = 863;
        test_data[1601] = 33'd3181973309;
        test_addr[1602] = 667;
        test_data[1602] = 33'd8159862793;
        test_addr[1603] = 668;
        test_data[1603] = 33'd4073128129;
        test_addr[1604] = 669;
        test_data[1604] = 33'd716422625;
        test_addr[1605] = 670;
        test_data[1605] = 33'd4276518473;
        test_addr[1606] = 671;
        test_data[1606] = 33'd2151985146;
        test_addr[1607] = 672;
        test_data[1607] = 33'd2838860096;
        test_addr[1608] = 673;
        test_data[1608] = 33'd2206060871;
        test_addr[1609] = 864;
        test_data[1609] = 33'd8417534796;
        test_addr[1610] = 865;
        test_data[1610] = 33'd2442557656;
        test_addr[1611] = 203;
        test_data[1611] = 33'd1831871360;
        test_addr[1612] = 866;
        test_data[1612] = 33'd2625374504;
        test_addr[1613] = 98;
        test_data[1613] = 33'd3514885588;
        test_addr[1614] = 99;
        test_data[1614] = 33'd3402368761;
        test_addr[1615] = 100;
        test_data[1615] = 33'd2034825318;
        test_addr[1616] = 101;
        test_data[1616] = 33'd4647523370;
        test_addr[1617] = 102;
        test_data[1617] = 33'd5031337076;
        test_addr[1618] = 103;
        test_data[1618] = 33'd437759945;
        test_addr[1619] = 104;
        test_data[1619] = 33'd3745214105;
        test_addr[1620] = 105;
        test_data[1620] = 33'd8171372023;
        test_addr[1621] = 106;
        test_data[1621] = 33'd4071584875;
        test_addr[1622] = 107;
        test_data[1622] = 33'd3862762663;
        test_addr[1623] = 108;
        test_data[1623] = 33'd7126178294;
        test_addr[1624] = 109;
        test_data[1624] = 33'd744992370;
        test_addr[1625] = 110;
        test_data[1625] = 33'd3882700174;
        test_addr[1626] = 111;
        test_data[1626] = 33'd1452439021;
        test_addr[1627] = 867;
        test_data[1627] = 33'd4191967086;
        test_addr[1628] = 868;
        test_data[1628] = 33'd5529877728;
        test_addr[1629] = 869;
        test_data[1629] = 33'd7275386462;
        test_addr[1630] = 870;
        test_data[1630] = 33'd5614271255;
        test_addr[1631] = 797;
        test_data[1631] = 33'd5823071774;
        test_addr[1632] = 798;
        test_data[1632] = 33'd4098353399;
        test_addr[1633] = 799;
        test_data[1633] = 33'd1518077955;
        test_addr[1634] = 800;
        test_data[1634] = 33'd754500382;
        test_addr[1635] = 801;
        test_data[1635] = 33'd8540563095;
        test_addr[1636] = 802;
        test_data[1636] = 33'd3063225216;
        test_addr[1637] = 803;
        test_data[1637] = 33'd1034772483;
        test_addr[1638] = 804;
        test_data[1638] = 33'd3999230770;
        test_addr[1639] = 805;
        test_data[1639] = 33'd2518139456;
        test_addr[1640] = 806;
        test_data[1640] = 33'd1466474561;
        test_addr[1641] = 807;
        test_data[1641] = 33'd639577463;
        test_addr[1642] = 808;
        test_data[1642] = 33'd4164035057;
        test_addr[1643] = 809;
        test_data[1643] = 33'd3968329823;
        test_addr[1644] = 810;
        test_data[1644] = 33'd8185367004;
        test_addr[1645] = 811;
        test_data[1645] = 33'd2968812544;
        test_addr[1646] = 812;
        test_data[1646] = 33'd2944629316;
        test_addr[1647] = 813;
        test_data[1647] = 33'd3207399348;
        test_addr[1648] = 814;
        test_data[1648] = 33'd2532614522;
        test_addr[1649] = 815;
        test_data[1649] = 33'd3596465989;
        test_addr[1650] = 816;
        test_data[1650] = 33'd2089907260;
        test_addr[1651] = 817;
        test_data[1651] = 33'd3539168386;
        test_addr[1652] = 818;
        test_data[1652] = 33'd6931281331;
        test_addr[1653] = 819;
        test_data[1653] = 33'd3407332409;
        test_addr[1654] = 820;
        test_data[1654] = 33'd4949092868;
        test_addr[1655] = 821;
        test_data[1655] = 33'd5071136119;
        test_addr[1656] = 822;
        test_data[1656] = 33'd4814794105;
        test_addr[1657] = 823;
        test_data[1657] = 33'd1941593249;
        test_addr[1658] = 824;
        test_data[1658] = 33'd4185437212;
        test_addr[1659] = 825;
        test_data[1659] = 33'd1444494147;
        test_addr[1660] = 826;
        test_data[1660] = 33'd293832577;
        test_addr[1661] = 827;
        test_data[1661] = 33'd4271161680;
        test_addr[1662] = 828;
        test_data[1662] = 33'd4228467133;
        test_addr[1663] = 829;
        test_data[1663] = 33'd2471067861;
        test_addr[1664] = 830;
        test_data[1664] = 33'd2151514164;
        test_addr[1665] = 871;
        test_data[1665] = 33'd8011412594;
        test_addr[1666] = 872;
        test_data[1666] = 33'd3833194746;
        test_addr[1667] = 482;
        test_data[1667] = 33'd3393357937;
        test_addr[1668] = 483;
        test_data[1668] = 33'd1323124837;
        test_addr[1669] = 484;
        test_data[1669] = 33'd998179708;
        test_addr[1670] = 485;
        test_data[1670] = 33'd1497784997;
        test_addr[1671] = 486;
        test_data[1671] = 33'd3551446877;
        test_addr[1672] = 487;
        test_data[1672] = 33'd4233924408;
        test_addr[1673] = 488;
        test_data[1673] = 33'd3230286556;
        test_addr[1674] = 489;
        test_data[1674] = 33'd654573334;
        test_addr[1675] = 490;
        test_data[1675] = 33'd7826218143;
        test_addr[1676] = 491;
        test_data[1676] = 33'd7857690380;
        test_addr[1677] = 492;
        test_data[1677] = 33'd2583156540;
        test_addr[1678] = 493;
        test_data[1678] = 33'd2880958133;
        test_addr[1679] = 494;
        test_data[1679] = 33'd1342614566;
        test_addr[1680] = 495;
        test_data[1680] = 33'd3753411143;
        test_addr[1681] = 496;
        test_data[1681] = 33'd3037540200;
        test_addr[1682] = 497;
        test_data[1682] = 33'd6905165754;
        test_addr[1683] = 498;
        test_data[1683] = 33'd4163492510;
        test_addr[1684] = 499;
        test_data[1684] = 33'd5671553493;
        test_addr[1685] = 500;
        test_data[1685] = 33'd1526412453;
        test_addr[1686] = 501;
        test_data[1686] = 33'd2592532499;
        test_addr[1687] = 502;
        test_data[1687] = 33'd1661402023;
        test_addr[1688] = 503;
        test_data[1688] = 33'd6034368094;
        test_addr[1689] = 504;
        test_data[1689] = 33'd225331988;
        test_addr[1690] = 873;
        test_data[1690] = 33'd5363552428;
        test_addr[1691] = 874;
        test_data[1691] = 33'd1199621947;
        test_addr[1692] = 875;
        test_data[1692] = 33'd2917729411;
        test_addr[1693] = 876;
        test_data[1693] = 33'd3736677355;
        test_addr[1694] = 877;
        test_data[1694] = 33'd6694736666;
        test_addr[1695] = 878;
        test_data[1695] = 33'd6221666340;
        test_addr[1696] = 879;
        test_data[1696] = 33'd4085858993;
        test_addr[1697] = 880;
        test_data[1697] = 33'd5402410262;
        test_addr[1698] = 881;
        test_data[1698] = 33'd3579846374;
        test_addr[1699] = 841;
        test_data[1699] = 33'd3495259579;
        test_addr[1700] = 842;
        test_data[1700] = 33'd1921393664;
        test_addr[1701] = 843;
        test_data[1701] = 33'd3444648562;
        test_addr[1702] = 882;
        test_data[1702] = 33'd386405139;
        test_addr[1703] = 883;
        test_data[1703] = 33'd1933304197;
        test_addr[1704] = 884;
        test_data[1704] = 33'd2315383485;
        test_addr[1705] = 885;
        test_data[1705] = 33'd3827515349;
        test_addr[1706] = 673;
        test_data[1706] = 33'd2206060871;
        test_addr[1707] = 674;
        test_data[1707] = 33'd5979601182;
        test_addr[1708] = 675;
        test_data[1708] = 33'd3430516374;
        test_addr[1709] = 676;
        test_data[1709] = 33'd662578081;
        test_addr[1710] = 677;
        test_data[1710] = 33'd6172600736;
        test_addr[1711] = 678;
        test_data[1711] = 33'd4202950769;
        test_addr[1712] = 679;
        test_data[1712] = 33'd6735495005;
        test_addr[1713] = 680;
        test_data[1713] = 33'd772379733;
        test_addr[1714] = 681;
        test_data[1714] = 33'd8296779550;
        test_addr[1715] = 886;
        test_data[1715] = 33'd4090995992;
        test_addr[1716] = 887;
        test_data[1716] = 33'd4779585778;
        test_addr[1717] = 888;
        test_data[1717] = 33'd1306365210;
        test_addr[1718] = 889;
        test_data[1718] = 33'd5823082263;
        test_addr[1719] = 890;
        test_data[1719] = 33'd5646568864;
        test_addr[1720] = 891;
        test_data[1720] = 33'd3155621446;
        test_addr[1721] = 892;
        test_data[1721] = 33'd5345881291;
        test_addr[1722] = 893;
        test_data[1722] = 33'd278268436;
        test_addr[1723] = 894;
        test_data[1723] = 33'd391382463;
        test_addr[1724] = 895;
        test_data[1724] = 33'd1907386417;
        test_addr[1725] = 896;
        test_data[1725] = 33'd1245387932;
        test_addr[1726] = 897;
        test_data[1726] = 33'd1758044350;
        test_addr[1727] = 898;
        test_data[1727] = 33'd8267258817;
        test_addr[1728] = 850;
        test_data[1728] = 33'd5039942209;
        test_addr[1729] = 851;
        test_data[1729] = 33'd7710705346;
        test_addr[1730] = 852;
        test_data[1730] = 33'd6999160267;
        test_addr[1731] = 853;
        test_data[1731] = 33'd8461085424;
        test_addr[1732] = 854;
        test_data[1732] = 33'd3331943895;
        test_addr[1733] = 855;
        test_data[1733] = 33'd1267612027;
        test_addr[1734] = 856;
        test_data[1734] = 33'd1996537634;
        test_addr[1735] = 857;
        test_data[1735] = 33'd4474236266;
        test_addr[1736] = 858;
        test_data[1736] = 33'd5019519486;
        test_addr[1737] = 859;
        test_data[1737] = 33'd3996213929;
        test_addr[1738] = 860;
        test_data[1738] = 33'd9740189;
        test_addr[1739] = 861;
        test_data[1739] = 33'd8539871332;
        test_addr[1740] = 862;
        test_data[1740] = 33'd8475427028;
        test_addr[1741] = 863;
        test_data[1741] = 33'd3181973309;
        test_addr[1742] = 864;
        test_data[1742] = 33'd4122567500;
        test_addr[1743] = 865;
        test_data[1743] = 33'd2442557656;
        test_addr[1744] = 866;
        test_data[1744] = 33'd4931277528;
        test_addr[1745] = 867;
        test_data[1745] = 33'd4191967086;
        test_addr[1746] = 899;
        test_data[1746] = 33'd6153803886;
        test_addr[1747] = 242;
        test_data[1747] = 33'd502196391;
        test_addr[1748] = 243;
        test_data[1748] = 33'd3483456815;
        test_addr[1749] = 244;
        test_data[1749] = 33'd1318439210;
        test_addr[1750] = 245;
        test_data[1750] = 33'd324506329;
        test_addr[1751] = 246;
        test_data[1751] = 33'd801919684;
        test_addr[1752] = 247;
        test_data[1752] = 33'd3793934249;
        test_addr[1753] = 248;
        test_data[1753] = 33'd5203023044;
        test_addr[1754] = 249;
        test_data[1754] = 33'd3317083412;
        test_addr[1755] = 250;
        test_data[1755] = 33'd1587295833;
        test_addr[1756] = 251;
        test_data[1756] = 33'd1245156121;
        test_addr[1757] = 252;
        test_data[1757] = 33'd855026393;
        test_addr[1758] = 253;
        test_data[1758] = 33'd2844318793;
        test_addr[1759] = 254;
        test_data[1759] = 33'd100893370;
        test_addr[1760] = 255;
        test_data[1760] = 33'd6802803139;
        test_addr[1761] = 256;
        test_data[1761] = 33'd2544636227;
        test_addr[1762] = 257;
        test_data[1762] = 33'd3530939413;
        test_addr[1763] = 258;
        test_data[1763] = 33'd5758805634;
        test_addr[1764] = 259;
        test_data[1764] = 33'd2333597655;
        test_addr[1765] = 260;
        test_data[1765] = 33'd1884041322;
        test_addr[1766] = 261;
        test_data[1766] = 33'd7353692545;
        test_addr[1767] = 262;
        test_data[1767] = 33'd3224676958;
        test_addr[1768] = 263;
        test_data[1768] = 33'd3200855956;
        test_addr[1769] = 264;
        test_data[1769] = 33'd4124826968;
        test_addr[1770] = 265;
        test_data[1770] = 33'd2848828629;
        test_addr[1771] = 266;
        test_data[1771] = 33'd2745001205;
        test_addr[1772] = 267;
        test_data[1772] = 33'd7924579505;
        test_addr[1773] = 900;
        test_data[1773] = 33'd3469687493;
        test_addr[1774] = 901;
        test_data[1774] = 33'd836715634;
        test_addr[1775] = 902;
        test_data[1775] = 33'd517865842;
        test_addr[1776] = 903;
        test_data[1776] = 33'd6825704132;
        test_addr[1777] = 904;
        test_data[1777] = 33'd3478950353;
        test_addr[1778] = 879;
        test_data[1778] = 33'd4085858993;
        test_addr[1779] = 880;
        test_data[1779] = 33'd1107442966;
        test_addr[1780] = 881;
        test_data[1780] = 33'd4979173725;
        test_addr[1781] = 882;
        test_data[1781] = 33'd6926039835;
        test_addr[1782] = 883;
        test_data[1782] = 33'd1933304197;
        test_addr[1783] = 884;
        test_data[1783] = 33'd2315383485;
        test_addr[1784] = 885;
        test_data[1784] = 33'd3827515349;
        test_addr[1785] = 886;
        test_data[1785] = 33'd4090995992;
        test_addr[1786] = 887;
        test_data[1786] = 33'd6066547373;
        test_addr[1787] = 888;
        test_data[1787] = 33'd1306365210;
        test_addr[1788] = 889;
        test_data[1788] = 33'd5311763766;
        test_addr[1789] = 890;
        test_data[1789] = 33'd1351601568;
        test_addr[1790] = 891;
        test_data[1790] = 33'd7338378116;
        test_addr[1791] = 892;
        test_data[1791] = 33'd1050913995;
        test_addr[1792] = 893;
        test_data[1792] = 33'd278268436;
        test_addr[1793] = 894;
        test_data[1793] = 33'd5600048239;
        test_addr[1794] = 895;
        test_data[1794] = 33'd4450168400;
        test_addr[1795] = 896;
        test_data[1795] = 33'd1245387932;
        test_addr[1796] = 897;
        test_data[1796] = 33'd8207417283;
        test_addr[1797] = 898;
        test_data[1797] = 33'd3972291521;
        test_addr[1798] = 899;
        test_data[1798] = 33'd1858836590;
        test_addr[1799] = 900;
        test_data[1799] = 33'd3469687493;
        test_addr[1800] = 905;
        test_data[1800] = 33'd4705211306;
        test_addr[1801] = 906;
        test_data[1801] = 33'd8513364149;
        test_addr[1802] = 907;
        test_data[1802] = 33'd6199781369;
        test_addr[1803] = 908;
        test_data[1803] = 33'd565450044;
        test_addr[1804] = 909;
        test_data[1804] = 33'd8570408910;
        test_addr[1805] = 910;
        test_data[1805] = 33'd1596033064;
        test_addr[1806] = 1004;
        test_data[1806] = 33'd2136110024;
        test_addr[1807] = 1005;
        test_data[1807] = 33'd2395804748;
        test_addr[1808] = 1006;
        test_data[1808] = 33'd479112565;
        test_addr[1809] = 1007;
        test_data[1809] = 33'd4059948122;
        test_addr[1810] = 1008;
        test_data[1810] = 33'd4049834946;
        test_addr[1811] = 1009;
        test_data[1811] = 33'd2905712961;
        test_addr[1812] = 1010;
        test_data[1812] = 33'd7097842582;
        test_addr[1813] = 1011;
        test_data[1813] = 33'd743506454;
        test_addr[1814] = 1012;
        test_data[1814] = 33'd891830012;
        test_addr[1815] = 1013;
        test_data[1815] = 33'd5345187767;
        test_addr[1816] = 1014;
        test_data[1816] = 33'd4755766292;
        test_addr[1817] = 1015;
        test_data[1817] = 33'd5963472566;
        test_addr[1818] = 1016;
        test_data[1818] = 33'd3935014123;
        test_addr[1819] = 1017;
        test_data[1819] = 33'd6325476189;
        test_addr[1820] = 1018;
        test_data[1820] = 33'd5064709768;
        test_addr[1821] = 1019;
        test_data[1821] = 33'd6033952536;
        test_addr[1822] = 1020;
        test_data[1822] = 33'd1804380535;
        test_addr[1823] = 1021;
        test_data[1823] = 33'd1888120797;
        test_addr[1824] = 1022;
        test_data[1824] = 33'd1248002737;
        test_addr[1825] = 1023;
        test_data[1825] = 33'd3621827067;
        test_addr[1826] = 0;
        test_data[1826] = 33'd3311723688;
        test_addr[1827] = 1;
        test_data[1827] = 33'd1830337710;
        test_addr[1828] = 2;
        test_data[1828] = 33'd2722018698;
        test_addr[1829] = 911;
        test_data[1829] = 33'd2521923331;
        test_addr[1830] = 912;
        test_data[1830] = 33'd3267133870;
        test_addr[1831] = 913;
        test_data[1831] = 33'd2193415700;
        test_addr[1832] = 914;
        test_data[1832] = 33'd284405744;
        test_addr[1833] = 915;
        test_data[1833] = 33'd839785297;
        test_addr[1834] = 916;
        test_data[1834] = 33'd3119093558;
        test_addr[1835] = 808;
        test_data[1835] = 33'd4164035057;
        test_addr[1836] = 809;
        test_data[1836] = 33'd3968329823;
        test_addr[1837] = 810;
        test_data[1837] = 33'd3890399708;
        test_addr[1838] = 811;
        test_data[1838] = 33'd2968812544;
        test_addr[1839] = 812;
        test_data[1839] = 33'd7027512201;
        test_addr[1840] = 813;
        test_data[1840] = 33'd3207399348;
        test_addr[1841] = 814;
        test_data[1841] = 33'd2532614522;
        test_addr[1842] = 815;
        test_data[1842] = 33'd3596465989;
        test_addr[1843] = 816;
        test_data[1843] = 33'd6554115366;
        test_addr[1844] = 817;
        test_data[1844] = 33'd3539168386;
        test_addr[1845] = 818;
        test_data[1845] = 33'd2636314035;
        test_addr[1846] = 917;
        test_data[1846] = 33'd8181607785;
        test_addr[1847] = 918;
        test_data[1847] = 33'd942389263;
        test_addr[1848] = 919;
        test_data[1848] = 33'd3709315097;
        test_addr[1849] = 920;
        test_data[1849] = 33'd8228993577;
        test_addr[1850] = 95;
        test_data[1850] = 33'd7638833046;
        test_addr[1851] = 96;
        test_data[1851] = 33'd6563312943;
        test_addr[1852] = 97;
        test_data[1852] = 33'd7961028460;
        test_addr[1853] = 98;
        test_data[1853] = 33'd8091935254;
        test_addr[1854] = 99;
        test_data[1854] = 33'd8113694733;
        test_addr[1855] = 100;
        test_data[1855] = 33'd2034825318;
        test_addr[1856] = 921;
        test_data[1856] = 33'd7347027749;
        test_addr[1857] = 922;
        test_data[1857] = 33'd6682095577;
        test_addr[1858] = 923;
        test_data[1858] = 33'd2212276299;
        test_addr[1859] = 924;
        test_data[1859] = 33'd7013976326;
        test_addr[1860] = 925;
        test_data[1860] = 33'd3444626246;
        test_addr[1861] = 926;
        test_data[1861] = 33'd8149379513;
        test_addr[1862] = 530;
        test_data[1862] = 33'd5401998960;
        test_addr[1863] = 531;
        test_data[1863] = 33'd1950799225;
        test_addr[1864] = 532;
        test_data[1864] = 33'd83719787;
        test_addr[1865] = 533;
        test_data[1865] = 33'd2895105766;
        test_addr[1866] = 534;
        test_data[1866] = 33'd2544290285;
        test_addr[1867] = 535;
        test_data[1867] = 33'd4594057720;
        test_addr[1868] = 536;
        test_data[1868] = 33'd2191918674;
        test_addr[1869] = 927;
        test_data[1869] = 33'd416978341;
        test_addr[1870] = 928;
        test_data[1870] = 33'd6743066105;
        test_addr[1871] = 929;
        test_data[1871] = 33'd3169898984;
        test_addr[1872] = 930;
        test_data[1872] = 33'd1164254761;
        test_addr[1873] = 931;
        test_data[1873] = 33'd4204922469;
        test_addr[1874] = 932;
        test_data[1874] = 33'd2044109763;
        test_addr[1875] = 933;
        test_data[1875] = 33'd3586314489;
        test_addr[1876] = 934;
        test_data[1876] = 33'd1840334227;
        test_addr[1877] = 935;
        test_data[1877] = 33'd2918620527;
        test_addr[1878] = 602;
        test_data[1878] = 33'd3640306504;
        test_addr[1879] = 603;
        test_data[1879] = 33'd2792617507;
        test_addr[1880] = 604;
        test_data[1880] = 33'd5293292067;
        test_addr[1881] = 605;
        test_data[1881] = 33'd1618144234;
        test_addr[1882] = 606;
        test_data[1882] = 33'd920782161;
        test_addr[1883] = 607;
        test_data[1883] = 33'd3986635328;
        test_addr[1884] = 608;
        test_data[1884] = 33'd2953791377;
        test_addr[1885] = 609;
        test_data[1885] = 33'd3511563354;
        test_addr[1886] = 610;
        test_data[1886] = 33'd2559326217;
        test_addr[1887] = 936;
        test_data[1887] = 33'd5501299366;
        test_addr[1888] = 937;
        test_data[1888] = 33'd1191377286;
        test_addr[1889] = 526;
        test_data[1889] = 33'd736640889;
        test_addr[1890] = 938;
        test_data[1890] = 33'd6638918666;
        test_addr[1891] = 939;
        test_data[1891] = 33'd775116840;
        test_addr[1892] = 940;
        test_data[1892] = 33'd8061157204;
        test_addr[1893] = 941;
        test_data[1893] = 33'd8527438570;
        test_addr[1894] = 942;
        test_data[1894] = 33'd5774807443;
        test_addr[1895] = 943;
        test_data[1895] = 33'd5172259901;
        test_addr[1896] = 944;
        test_data[1896] = 33'd4223266270;
        test_addr[1897] = 945;
        test_data[1897] = 33'd2788157755;
        test_addr[1898] = 946;
        test_data[1898] = 33'd2141896945;
        test_addr[1899] = 947;
        test_data[1899] = 33'd7419450515;
        test_addr[1900] = 948;
        test_data[1900] = 33'd1116008264;
        test_addr[1901] = 949;
        test_data[1901] = 33'd4425696288;
        test_addr[1902] = 950;
        test_data[1902] = 33'd2097728883;
        test_addr[1903] = 951;
        test_data[1903] = 33'd5511087095;
        test_addr[1904] = 952;
        test_data[1904] = 33'd1618745728;
        test_addr[1905] = 953;
        test_data[1905] = 33'd8202780824;
        test_addr[1906] = 954;
        test_data[1906] = 33'd3692314337;
        test_addr[1907] = 955;
        test_data[1907] = 33'd6120939512;
        test_addr[1908] = 956;
        test_data[1908] = 33'd2529817444;
        test_addr[1909] = 957;
        test_data[1909] = 33'd2432425057;
        test_addr[1910] = 958;
        test_data[1910] = 33'd5731383527;
        test_addr[1911] = 959;
        test_data[1911] = 33'd1670570220;
        test_addr[1912] = 453;
        test_data[1912] = 33'd4144249236;
        test_addr[1913] = 454;
        test_data[1913] = 33'd3006483553;
        test_addr[1914] = 455;
        test_data[1914] = 33'd3480902115;
        test_addr[1915] = 456;
        test_data[1915] = 33'd6689270127;
        test_addr[1916] = 457;
        test_data[1916] = 33'd7177631868;
        test_addr[1917] = 960;
        test_data[1917] = 33'd269126776;
        test_addr[1918] = 793;
        test_data[1918] = 33'd8088053104;
        test_addr[1919] = 794;
        test_data[1919] = 33'd4491353472;
        test_addr[1920] = 795;
        test_data[1920] = 33'd2128607902;
        test_addr[1921] = 796;
        test_data[1921] = 33'd4275211649;
        test_addr[1922] = 797;
        test_data[1922] = 33'd1528104478;
        test_addr[1923] = 798;
        test_data[1923] = 33'd4098353399;
        test_addr[1924] = 799;
        test_data[1924] = 33'd1518077955;
        test_addr[1925] = 800;
        test_data[1925] = 33'd4949084106;
        test_addr[1926] = 801;
        test_data[1926] = 33'd6140785602;
        test_addr[1927] = 961;
        test_data[1927] = 33'd1162456992;
        test_addr[1928] = 962;
        test_data[1928] = 33'd7258591980;
        test_addr[1929] = 963;
        test_data[1929] = 33'd3714607084;
        test_addr[1930] = 964;
        test_data[1930] = 33'd2358691;
        test_addr[1931] = 965;
        test_data[1931] = 33'd3011036640;
        test_addr[1932] = 333;
        test_data[1932] = 33'd2296982685;
        test_addr[1933] = 334;
        test_data[1933] = 33'd6237591288;
        test_addr[1934] = 335;
        test_data[1934] = 33'd1195626943;
        test_addr[1935] = 336;
        test_data[1935] = 33'd1688024943;
        test_addr[1936] = 337;
        test_data[1936] = 33'd750261429;
        test_addr[1937] = 338;
        test_data[1937] = 33'd1821314294;
        test_addr[1938] = 339;
        test_data[1938] = 33'd8261343235;
        test_addr[1939] = 340;
        test_data[1939] = 33'd1638179589;
        test_addr[1940] = 341;
        test_data[1940] = 33'd315843574;
        test_addr[1941] = 342;
        test_data[1941] = 33'd4716402424;
        test_addr[1942] = 343;
        test_data[1942] = 33'd2846218665;
        test_addr[1943] = 344;
        test_data[1943] = 33'd768223443;
        test_addr[1944] = 345;
        test_data[1944] = 33'd2791959723;
        test_addr[1945] = 346;
        test_data[1945] = 33'd3770003965;
        test_addr[1946] = 347;
        test_data[1946] = 33'd4150740891;
        test_addr[1947] = 348;
        test_data[1947] = 33'd904943400;
        test_addr[1948] = 349;
        test_data[1948] = 33'd8458599857;
        test_addr[1949] = 350;
        test_data[1949] = 33'd617222912;
        test_addr[1950] = 351;
        test_data[1950] = 33'd7647554633;
        test_addr[1951] = 352;
        test_data[1951] = 33'd163922335;
        test_addr[1952] = 353;
        test_data[1952] = 33'd8435705399;
        test_addr[1953] = 354;
        test_data[1953] = 33'd4080977870;
        test_addr[1954] = 355;
        test_data[1954] = 33'd7454752690;
        test_addr[1955] = 356;
        test_data[1955] = 33'd2257235136;
        test_addr[1956] = 357;
        test_data[1956] = 33'd8410799578;
        test_addr[1957] = 358;
        test_data[1957] = 33'd3685422029;
        test_addr[1958] = 359;
        test_data[1958] = 33'd8202096931;
        test_addr[1959] = 360;
        test_data[1959] = 33'd4497849208;
        test_addr[1960] = 361;
        test_data[1960] = 33'd2414551097;
        test_addr[1961] = 362;
        test_data[1961] = 33'd5289004044;
        test_addr[1962] = 363;
        test_data[1962] = 33'd2723076636;
        test_addr[1963] = 364;
        test_data[1963] = 33'd1333182938;
        test_addr[1964] = 966;
        test_data[1964] = 33'd2186720106;
        test_addr[1965] = 967;
        test_data[1965] = 33'd6957448563;
        test_addr[1966] = 968;
        test_data[1966] = 33'd8031544118;
        test_addr[1967] = 969;
        test_data[1967] = 33'd3579876324;
        test_addr[1968] = 970;
        test_data[1968] = 33'd2846411311;
        test_addr[1969] = 971;
        test_data[1969] = 33'd3021945945;
        test_addr[1970] = 972;
        test_data[1970] = 33'd7446923207;
        test_addr[1971] = 973;
        test_data[1971] = 33'd6606993614;
        test_addr[1972] = 974;
        test_data[1972] = 33'd2563567935;
        test_addr[1973] = 975;
        test_data[1973] = 33'd267738865;
        test_addr[1974] = 976;
        test_data[1974] = 33'd5063658287;
        test_addr[1975] = 977;
        test_data[1975] = 33'd380731391;
        test_addr[1976] = 978;
        test_data[1976] = 33'd2323391226;
        test_addr[1977] = 979;
        test_data[1977] = 33'd3960867072;
        test_addr[1978] = 980;
        test_data[1978] = 33'd6929535015;
        test_addr[1979] = 981;
        test_data[1979] = 33'd2623441966;
        test_addr[1980] = 982;
        test_data[1980] = 33'd8533471868;
        test_addr[1981] = 983;
        test_data[1981] = 33'd3660155862;
        test_addr[1982] = 458;
        test_data[1982] = 33'd4143306261;
        test_addr[1983] = 459;
        test_data[1983] = 33'd1894780540;
        test_addr[1984] = 460;
        test_data[1984] = 33'd2715526497;
        test_addr[1985] = 461;
        test_data[1985] = 33'd2207510278;
        test_addr[1986] = 462;
        test_data[1986] = 33'd2318869365;
        test_addr[1987] = 463;
        test_data[1987] = 33'd909928079;
        test_addr[1988] = 464;
        test_data[1988] = 33'd3521762258;
        test_addr[1989] = 465;
        test_data[1989] = 33'd4173322230;
        test_addr[1990] = 466;
        test_data[1990] = 33'd1591617322;
        test_addr[1991] = 467;
        test_data[1991] = 33'd5257053311;
        test_addr[1992] = 984;
        test_data[1992] = 33'd978931367;
        test_addr[1993] = 985;
        test_data[1993] = 33'd957211627;
        test_addr[1994] = 115;
        test_data[1994] = 33'd1652892941;
        test_addr[1995] = 116;
        test_data[1995] = 33'd6669989840;
        test_addr[1996] = 117;
        test_data[1996] = 33'd4220214550;
        test_addr[1997] = 118;
        test_data[1997] = 33'd852272656;
        test_addr[1998] = 119;
        test_data[1998] = 33'd4958189913;
        test_addr[1999] = 120;
        test_data[1999] = 33'd5122421660;
        test_addr[2000] = 121;
        test_data[2000] = 33'd2605200182;
        test_addr[2001] = 986;
        test_data[2001] = 33'd3822672388;
        test_addr[2002] = 987;
        test_data[2002] = 33'd7830660222;
        test_addr[2003] = 342;
        test_data[2003] = 33'd421435128;
        test_addr[2004] = 343;
        test_data[2004] = 33'd2846218665;
        test_addr[2005] = 344;
        test_data[2005] = 33'd768223443;
        test_addr[2006] = 345;
        test_data[2006] = 33'd2791959723;
        test_addr[2007] = 346;
        test_data[2007] = 33'd3770003965;
        test_addr[2008] = 347;
        test_data[2008] = 33'd4150740891;
        test_addr[2009] = 348;
        test_data[2009] = 33'd904943400;
        test_addr[2010] = 349;
        test_data[2010] = 33'd4163632561;
        test_addr[2011] = 350;
        test_data[2011] = 33'd617222912;
        test_addr[2012] = 351;
        test_data[2012] = 33'd5000043653;
        test_addr[2013] = 352;
        test_data[2013] = 33'd163922335;
        test_addr[2014] = 353;
        test_data[2014] = 33'd7285498847;
        test_addr[2015] = 354;
        test_data[2015] = 33'd4080977870;
        test_addr[2016] = 355;
        test_data[2016] = 33'd7270526247;
        test_addr[2017] = 356;
        test_data[2017] = 33'd2257235136;
        test_addr[2018] = 357;
        test_data[2018] = 33'd4115832282;
        test_addr[2019] = 358;
        test_data[2019] = 33'd3685422029;
        test_addr[2020] = 359;
        test_data[2020] = 33'd3907129635;
        test_addr[2021] = 360;
        test_data[2021] = 33'd202881912;
        test_addr[2022] = 361;
        test_data[2022] = 33'd2414551097;
        test_addr[2023] = 362;
        test_data[2023] = 33'd4372899909;
        test_addr[2024] = 988;
        test_data[2024] = 33'd3995363066;
        test_addr[2025] = 989;
        test_data[2025] = 33'd4181739735;
        test_addr[2026] = 990;
        test_data[2026] = 33'd6827955185;
        test_addr[2027] = 991;
        test_data[2027] = 33'd88478458;
        test_addr[2028] = 992;
        test_data[2028] = 33'd669592020;
        test_addr[2029] = 993;
        test_data[2029] = 33'd1916779651;
        test_addr[2030] = 994;
        test_data[2030] = 33'd7204141108;
        test_addr[2031] = 196;
        test_data[2031] = 33'd2584950764;
        test_addr[2032] = 197;
        test_data[2032] = 33'd1696743885;
        test_addr[2033] = 198;
        test_data[2033] = 33'd2875093575;
        test_addr[2034] = 199;
        test_data[2034] = 33'd117868309;
        test_addr[2035] = 200;
        test_data[2035] = 33'd4066794897;
        test_addr[2036] = 201;
        test_data[2036] = 33'd5774316157;
        test_addr[2037] = 202;
        test_data[2037] = 33'd1056869093;
        test_addr[2038] = 995;
        test_data[2038] = 33'd55503118;
        test_addr[2039] = 996;
        test_data[2039] = 33'd1855610634;
        test_addr[2040] = 997;
        test_data[2040] = 33'd2243105101;
        test_addr[2041] = 998;
        test_data[2041] = 33'd8470231622;
        test_addr[2042] = 999;
        test_data[2042] = 33'd1429796383;
        test_addr[2043] = 1000;
        test_data[2043] = 33'd136122382;
        test_addr[2044] = 1001;
        test_data[2044] = 33'd1757685921;
        test_addr[2045] = 1002;
        test_data[2045] = 33'd1476013580;
        test_addr[2046] = 1003;
        test_data[2046] = 33'd1864759393;
        test_addr[2047] = 1004;
        test_data[2047] = 33'd7493196472;
        test_addr[2048] = 1005;
        test_data[2048] = 33'd2395804748;
        test_addr[2049] = 1006;
        test_data[2049] = 33'd479112565;
        test_addr[2050] = 1007;
        test_data[2050] = 33'd4059948122;
        test_addr[2051] = 1008;
        test_data[2051] = 33'd4049834946;
        test_addr[2052] = 1009;
        test_data[2052] = 33'd2905712961;
        test_addr[2053] = 86;
        test_data[2053] = 33'd5256286182;
        test_addr[2054] = 87;
        test_data[2054] = 33'd1074381877;
        test_addr[2055] = 88;
        test_data[2055] = 33'd1562271896;
        test_addr[2056] = 1010;
        test_data[2056] = 33'd4496809828;
        test_addr[2057] = 1011;
        test_data[2057] = 33'd743506454;
        test_addr[2058] = 1012;
        test_data[2058] = 33'd891830012;
        test_addr[2059] = 686;
        test_data[2059] = 33'd4109187007;
        test_addr[2060] = 1013;
        test_data[2060] = 33'd1050220471;
        test_addr[2061] = 517;
        test_data[2061] = 33'd6337423047;
        test_addr[2062] = 518;
        test_data[2062] = 33'd849664853;
        test_addr[2063] = 519;
        test_data[2063] = 33'd4049498241;
        test_addr[2064] = 520;
        test_data[2064] = 33'd7289269808;
        test_addr[2065] = 521;
        test_data[2065] = 33'd3220870596;
        test_addr[2066] = 522;
        test_data[2066] = 33'd3048636483;
        test_addr[2067] = 523;
        test_data[2067] = 33'd1382851467;
        test_addr[2068] = 524;
        test_data[2068] = 33'd8075586282;
        test_addr[2069] = 525;
        test_data[2069] = 33'd2281015751;
        test_addr[2070] = 526;
        test_data[2070] = 33'd736640889;
        test_addr[2071] = 527;
        test_data[2071] = 33'd3884199812;
        test_addr[2072] = 528;
        test_data[2072] = 33'd2463388950;
        test_addr[2073] = 529;
        test_data[2073] = 33'd4484867377;
        test_addr[2074] = 530;
        test_data[2074] = 33'd1107031664;
        test_addr[2075] = 531;
        test_data[2075] = 33'd1950799225;
        test_addr[2076] = 532;
        test_data[2076] = 33'd83719787;
        test_addr[2077] = 533;
        test_data[2077] = 33'd2895105766;
        test_addr[2078] = 534;
        test_data[2078] = 33'd6961196210;
        test_addr[2079] = 535;
        test_data[2079] = 33'd7081777176;
        test_addr[2080] = 536;
        test_data[2080] = 33'd5274069176;
        test_addr[2081] = 537;
        test_data[2081] = 33'd1269482248;
        test_addr[2082] = 538;
        test_data[2082] = 33'd2662158238;
        test_addr[2083] = 1014;
        test_data[2083] = 33'd460798996;
        test_addr[2084] = 1015;
        test_data[2084] = 33'd1668505270;
        test_addr[2085] = 916;
        test_data[2085] = 33'd3119093558;
        test_addr[2086] = 917;
        test_data[2086] = 33'd3886640489;
        test_addr[2087] = 918;
        test_data[2087] = 33'd5066764034;
        test_addr[2088] = 919;
        test_data[2088] = 33'd3709315097;
        test_addr[2089] = 920;
        test_data[2089] = 33'd3934026281;
        test_addr[2090] = 921;
        test_data[2090] = 33'd3052060453;
        test_addr[2091] = 922;
        test_data[2091] = 33'd2387128281;
        test_addr[2092] = 923;
        test_data[2092] = 33'd2212276299;
        test_addr[2093] = 924;
        test_data[2093] = 33'd6610014572;
        test_addr[2094] = 925;
        test_data[2094] = 33'd3444626246;
        test_addr[2095] = 926;
        test_data[2095] = 33'd5812108424;
        test_addr[2096] = 927;
        test_data[2096] = 33'd4446365110;
        test_addr[2097] = 928;
        test_data[2097] = 33'd2448098809;
        test_addr[2098] = 929;
        test_data[2098] = 33'd3169898984;
        test_addr[2099] = 930;
        test_data[2099] = 33'd4474769448;
        test_addr[2100] = 931;
        test_data[2100] = 33'd4341127265;
        test_addr[2101] = 932;
        test_data[2101] = 33'd5265225828;
        test_addr[2102] = 933;
        test_data[2102] = 33'd8484648228;
        test_addr[2103] = 934;
        test_data[2103] = 33'd1840334227;
        test_addr[2104] = 935;
        test_data[2104] = 33'd2918620527;
        test_addr[2105] = 936;
        test_data[2105] = 33'd1206332070;
        test_addr[2106] = 937;
        test_data[2106] = 33'd1191377286;
        test_addr[2107] = 938;
        test_data[2107] = 33'd8199942467;
        test_addr[2108] = 939;
        test_data[2108] = 33'd775116840;
        test_addr[2109] = 940;
        test_data[2109] = 33'd3766189908;
        test_addr[2110] = 941;
        test_data[2110] = 33'd4232471274;
        test_addr[2111] = 942;
        test_data[2111] = 33'd1479840147;
        test_addr[2112] = 943;
        test_data[2112] = 33'd877292605;
        test_addr[2113] = 944;
        test_data[2113] = 33'd4223266270;
        test_addr[2114] = 945;
        test_data[2114] = 33'd2788157755;
        test_addr[2115] = 946;
        test_data[2115] = 33'd5634699405;
        test_addr[2116] = 947;
        test_data[2116] = 33'd3124483219;
        test_addr[2117] = 948;
        test_data[2117] = 33'd1116008264;
        test_addr[2118] = 949;
        test_data[2118] = 33'd5432910093;
        test_addr[2119] = 950;
        test_data[2119] = 33'd8309881675;
        test_addr[2120] = 951;
        test_data[2120] = 33'd1216119799;
        test_addr[2121] = 952;
        test_data[2121] = 33'd4376601232;
        test_addr[2122] = 953;
        test_data[2122] = 33'd3907813528;
        test_addr[2123] = 954;
        test_data[2123] = 33'd3692314337;
        test_addr[2124] = 955;
        test_data[2124] = 33'd1825972216;
        test_addr[2125] = 1016;
        test_data[2125] = 33'd7356750345;
        test_addr[2126] = 1017;
        test_data[2126] = 33'd4588675422;
        test_addr[2127] = 1018;
        test_data[2127] = 33'd4561150164;
        test_addr[2128] = 1019;
        test_data[2128] = 33'd1738985240;
        test_addr[2129] = 664;
        test_data[2129] = 33'd4123313617;
        test_addr[2130] = 665;
        test_data[2130] = 33'd1234201857;
        test_addr[2131] = 666;
        test_data[2131] = 33'd4740404902;
        test_addr[2132] = 667;
        test_data[2132] = 33'd5799315301;
        test_addr[2133] = 668;
        test_data[2133] = 33'd7628276364;
        test_addr[2134] = 669;
        test_data[2134] = 33'd716422625;
        test_addr[2135] = 670;
        test_data[2135] = 33'd4276518473;
        test_addr[2136] = 671;
        test_data[2136] = 33'd7126837724;
        test_addr[2137] = 672;
        test_data[2137] = 33'd2838860096;
        test_addr[2138] = 673;
        test_data[2138] = 33'd2206060871;
        test_addr[2139] = 674;
        test_data[2139] = 33'd1684633886;
        test_addr[2140] = 675;
        test_data[2140] = 33'd7789829779;
        test_addr[2141] = 676;
        test_data[2141] = 33'd662578081;
        test_addr[2142] = 677;
        test_data[2142] = 33'd1877633440;
        test_addr[2143] = 678;
        test_data[2143] = 33'd4202950769;
        test_addr[2144] = 679;
        test_data[2144] = 33'd6532134520;
        test_addr[2145] = 680;
        test_data[2145] = 33'd772379733;
        test_addr[2146] = 681;
        test_data[2146] = 33'd7492785302;
        test_addr[2147] = 682;
        test_data[2147] = 33'd666405120;
        test_addr[2148] = 683;
        test_data[2148] = 33'd1731237928;
        test_addr[2149] = 684;
        test_data[2149] = 33'd7720316730;
        test_addr[2150] = 685;
        test_data[2150] = 33'd4766112059;
        test_addr[2151] = 686;
        test_data[2151] = 33'd4109187007;
        test_addr[2152] = 687;
        test_data[2152] = 33'd7538684182;
        test_addr[2153] = 688;
        test_data[2153] = 33'd2293783707;
        test_addr[2154] = 689;
        test_data[2154] = 33'd5422559078;
        test_addr[2155] = 690;
        test_data[2155] = 33'd96841274;
        test_addr[2156] = 691;
        test_data[2156] = 33'd3289493552;
        test_addr[2157] = 692;
        test_data[2157] = 33'd4364113395;
        test_addr[2158] = 693;
        test_data[2158] = 33'd2076034828;
        test_addr[2159] = 1020;
        test_data[2159] = 33'd1804380535;
        test_addr[2160] = 1021;
        test_data[2160] = 33'd1888120797;
        test_addr[2161] = 1022;
        test_data[2161] = 33'd1248002737;
        test_addr[2162] = 1023;
        test_data[2162] = 33'd7969163955;
        test_addr[2163] = 0;
        test_data[2163] = 33'd3311723688;
        test_addr[2164] = 1;
        test_data[2164] = 33'd1830337710;
        test_addr[2165] = 2;
        test_data[2165] = 33'd5023780917;
        test_addr[2166] = 3;
        test_data[2166] = 33'd2095642455;
        test_addr[2167] = 4;
        test_data[2167] = 33'd5220581012;
        test_addr[2168] = 5;
        test_data[2168] = 33'd4780945538;
        test_addr[2169] = 6;
        test_data[2169] = 33'd3199283968;
        test_addr[2170] = 7;
        test_data[2170] = 33'd966600747;
        test_addr[2171] = 8;
        test_data[2171] = 33'd7673366633;
        test_addr[2172] = 9;
        test_data[2172] = 33'd6432748424;
        test_addr[2173] = 10;
        test_data[2173] = 33'd2701436524;
        test_addr[2174] = 11;
        test_data[2174] = 33'd142496755;
        test_addr[2175] = 12;
        test_data[2175] = 33'd1442523325;
        test_addr[2176] = 834;
        test_data[2176] = 33'd1624961981;
        test_addr[2177] = 835;
        test_data[2177] = 33'd7328249927;
        test_addr[2178] = 836;
        test_data[2178] = 33'd7783696041;
        test_addr[2179] = 837;
        test_data[2179] = 33'd2295011618;
        test_addr[2180] = 838;
        test_data[2180] = 33'd2598268969;
        test_addr[2181] = 839;
        test_data[2181] = 33'd6692521765;
        test_addr[2182] = 840;
        test_data[2182] = 33'd2690967453;
        test_addr[2183] = 841;
        test_data[2183] = 33'd3495259579;
        test_addr[2184] = 842;
        test_data[2184] = 33'd7924678908;
        test_addr[2185] = 843;
        test_data[2185] = 33'd3444648562;
        test_addr[2186] = 844;
        test_data[2186] = 33'd5728272940;
        test_addr[2187] = 13;
        test_data[2187] = 33'd2440374455;
        test_addr[2188] = 14;
        test_data[2188] = 33'd1328303385;
        test_addr[2189] = 15;
        test_data[2189] = 33'd8149460789;
        test_addr[2190] = 16;
        test_data[2190] = 33'd38352283;
        test_addr[2191] = 17;
        test_data[2191] = 33'd332043326;
        test_addr[2192] = 18;
        test_data[2192] = 33'd6967006121;
        test_addr[2193] = 19;
        test_data[2193] = 33'd3066389384;
        test_addr[2194] = 406;
        test_data[2194] = 33'd8565236662;
        test_addr[2195] = 407;
        test_data[2195] = 33'd3650981421;
        test_addr[2196] = 408;
        test_data[2196] = 33'd1991242564;
        test_addr[2197] = 409;
        test_data[2197] = 33'd881702054;
        test_addr[2198] = 410;
        test_data[2198] = 33'd3442998655;
        test_addr[2199] = 411;
        test_data[2199] = 33'd5670175044;
        test_addr[2200] = 412;
        test_data[2200] = 33'd3063633923;
        test_addr[2201] = 413;
        test_data[2201] = 33'd6853723507;
        test_addr[2202] = 414;
        test_data[2202] = 33'd2622463751;
        test_addr[2203] = 20;
        test_data[2203] = 33'd2016265322;
        test_addr[2204] = 848;
        test_data[2204] = 33'd2055262394;
        test_addr[2205] = 849;
        test_data[2205] = 33'd8383173157;
        test_addr[2206] = 850;
        test_data[2206] = 33'd7945378706;
        test_addr[2207] = 851;
        test_data[2207] = 33'd3415738050;
        test_addr[2208] = 852;
        test_data[2208] = 33'd2704192971;
        test_addr[2209] = 853;
        test_data[2209] = 33'd5362019442;
        test_addr[2210] = 854;
        test_data[2210] = 33'd3331943895;
        test_addr[2211] = 855;
        test_data[2211] = 33'd1267612027;
        test_addr[2212] = 856;
        test_data[2212] = 33'd5116504764;
        test_addr[2213] = 21;
        test_data[2213] = 33'd2004948545;
        test_addr[2214] = 22;
        test_data[2214] = 33'd7944965326;
        test_addr[2215] = 23;
        test_data[2215] = 33'd36425900;
        test_addr[2216] = 595;
        test_data[2216] = 33'd5529106125;
        test_addr[2217] = 596;
        test_data[2217] = 33'd1972695031;
        test_addr[2218] = 597;
        test_data[2218] = 33'd3535940700;
        test_addr[2219] = 598;
        test_data[2219] = 33'd4111524620;
        test_addr[2220] = 599;
        test_data[2220] = 33'd6471392202;
        test_addr[2221] = 600;
        test_data[2221] = 33'd3084518942;
        test_addr[2222] = 601;
        test_data[2222] = 33'd1061024359;
        test_addr[2223] = 602;
        test_data[2223] = 33'd8519798258;
        test_addr[2224] = 603;
        test_data[2224] = 33'd2792617507;
        test_addr[2225] = 24;
        test_data[2225] = 33'd759408867;
        test_addr[2226] = 25;
        test_data[2226] = 33'd2632895408;
        test_addr[2227] = 316;
        test_data[2227] = 33'd8408132505;
        test_addr[2228] = 317;
        test_data[2228] = 33'd2374556068;
        test_addr[2229] = 318;
        test_data[2229] = 33'd5960843327;
        test_addr[2230] = 319;
        test_data[2230] = 33'd357113237;
        test_addr[2231] = 320;
        test_data[2231] = 33'd2364460379;
        test_addr[2232] = 321;
        test_data[2232] = 33'd4278979725;
        test_addr[2233] = 322;
        test_data[2233] = 33'd341336502;
        test_addr[2234] = 323;
        test_data[2234] = 33'd1953799233;
        test_addr[2235] = 26;
        test_data[2235] = 33'd3295931461;
        test_addr[2236] = 408;
        test_data[2236] = 33'd1991242564;
        test_addr[2237] = 409;
        test_data[2237] = 33'd881702054;
        test_addr[2238] = 410;
        test_data[2238] = 33'd3442998655;
        test_addr[2239] = 27;
        test_data[2239] = 33'd5174133089;
        test_addr[2240] = 28;
        test_data[2240] = 33'd4574886892;
        test_addr[2241] = 29;
        test_data[2241] = 33'd7841180695;
        test_addr[2242] = 30;
        test_data[2242] = 33'd3059136363;
        test_addr[2243] = 31;
        test_data[2243] = 33'd1175891688;
        test_addr[2244] = 32;
        test_data[2244] = 33'd8171421984;
        test_addr[2245] = 33;
        test_data[2245] = 33'd6087571875;
        test_addr[2246] = 34;
        test_data[2246] = 33'd5764074333;
        test_addr[2247] = 35;
        test_data[2247] = 33'd5855191057;
        test_addr[2248] = 36;
        test_data[2248] = 33'd4012222965;
        test_addr[2249] = 37;
        test_data[2249] = 33'd6469038085;
        test_addr[2250] = 38;
        test_data[2250] = 33'd203837415;
        test_addr[2251] = 39;
        test_data[2251] = 33'd4702211103;
        test_addr[2252] = 40;
        test_data[2252] = 33'd5826054394;
        test_addr[2253] = 41;
        test_data[2253] = 33'd7578358043;
        test_addr[2254] = 42;
        test_data[2254] = 33'd3684409809;
        test_addr[2255] = 43;
        test_data[2255] = 33'd2514013501;
        test_addr[2256] = 44;
        test_data[2256] = 33'd3264450694;
        test_addr[2257] = 45;
        test_data[2257] = 33'd124332228;
        test_addr[2258] = 46;
        test_data[2258] = 33'd733918119;
        test_addr[2259] = 47;
        test_data[2259] = 33'd2276482309;
        test_addr[2260] = 48;
        test_data[2260] = 33'd6922508808;
        test_addr[2261] = 49;
        test_data[2261] = 33'd3795521150;
        test_addr[2262] = 50;
        test_data[2262] = 33'd6975386861;
        test_addr[2263] = 51;
        test_data[2263] = 33'd3965955358;
        test_addr[2264] = 52;
        test_data[2264] = 33'd7687114890;
        test_addr[2265] = 53;
        test_data[2265] = 33'd1370932658;
        test_addr[2266] = 54;
        test_data[2266] = 33'd3762196439;
        test_addr[2267] = 55;
        test_data[2267] = 33'd3541808763;
        test_addr[2268] = 56;
        test_data[2268] = 33'd6823173999;
        test_addr[2269] = 57;
        test_data[2269] = 33'd3015078990;
        test_addr[2270] = 58;
        test_data[2270] = 33'd7633147289;
        test_addr[2271] = 59;
        test_data[2271] = 33'd8267524516;
        test_addr[2272] = 60;
        test_data[2272] = 33'd2524153113;
        test_addr[2273] = 61;
        test_data[2273] = 33'd2579925800;
        test_addr[2274] = 62;
        test_data[2274] = 33'd6096172882;
        test_addr[2275] = 63;
        test_data[2275] = 33'd1646915880;
        test_addr[2276] = 64;
        test_data[2276] = 33'd1966218068;
        test_addr[2277] = 665;
        test_data[2277] = 33'd1234201857;
        test_addr[2278] = 666;
        test_data[2278] = 33'd4733086078;
        test_addr[2279] = 65;
        test_data[2279] = 33'd1845517365;
        test_addr[2280] = 66;
        test_data[2280] = 33'd2814571527;
        test_addr[2281] = 67;
        test_data[2281] = 33'd6291224010;
        test_addr[2282] = 68;
        test_data[2282] = 33'd4069819184;
        test_addr[2283] = 69;
        test_data[2283] = 33'd4483095371;
        test_addr[2284] = 70;
        test_data[2284] = 33'd2049921272;
        test_addr[2285] = 71;
        test_data[2285] = 33'd7707500985;
        test_addr[2286] = 72;
        test_data[2286] = 33'd1234549181;
        test_addr[2287] = 73;
        test_data[2287] = 33'd8377247341;
        test_addr[2288] = 74;
        test_data[2288] = 33'd4823463627;
        test_addr[2289] = 75;
        test_data[2289] = 33'd5407702443;
        test_addr[2290] = 76;
        test_data[2290] = 33'd1083302262;
        test_addr[2291] = 77;
        test_data[2291] = 33'd2876543838;
        test_addr[2292] = 78;
        test_data[2292] = 33'd3671955214;
        test_addr[2293] = 79;
        test_data[2293] = 33'd238733017;
        test_addr[2294] = 80;
        test_data[2294] = 33'd2907114715;
        test_addr[2295] = 81;
        test_data[2295] = 33'd1759133022;
        test_addr[2296] = 82;
        test_data[2296] = 33'd2394041630;
        test_addr[2297] = 83;
        test_data[2297] = 33'd2532816163;
        test_addr[2298] = 84;
        test_data[2298] = 33'd655204540;
        test_addr[2299] = 85;
        test_data[2299] = 33'd4108519334;
        test_addr[2300] = 86;
        test_data[2300] = 33'd6178761991;
        test_addr[2301] = 214;
        test_data[2301] = 33'd635033231;
        test_addr[2302] = 215;
        test_data[2302] = 33'd4098659685;
        test_addr[2303] = 216;
        test_data[2303] = 33'd1581642574;
        test_addr[2304] = 217;
        test_data[2304] = 33'd2718828492;
        test_addr[2305] = 218;
        test_data[2305] = 33'd1056999408;
        test_addr[2306] = 219;
        test_data[2306] = 33'd5813290370;
        test_addr[2307] = 220;
        test_data[2307] = 33'd5067496498;
        test_addr[2308] = 221;
        test_data[2308] = 33'd3019464660;
        test_addr[2309] = 222;
        test_data[2309] = 33'd1384897455;
        test_addr[2310] = 223;
        test_data[2310] = 33'd1381153484;
        test_addr[2311] = 224;
        test_data[2311] = 33'd463140193;
        test_addr[2312] = 225;
        test_data[2312] = 33'd1457651049;
        test_addr[2313] = 226;
        test_data[2313] = 33'd7610345369;
        test_addr[2314] = 227;
        test_data[2314] = 33'd2688484918;
        test_addr[2315] = 228;
        test_data[2315] = 33'd4120475529;
        test_addr[2316] = 229;
        test_data[2316] = 33'd665005425;
        test_addr[2317] = 230;
        test_data[2317] = 33'd988458485;
        test_addr[2318] = 231;
        test_data[2318] = 33'd6165527530;
        test_addr[2319] = 232;
        test_data[2319] = 33'd1665029119;
        test_addr[2320] = 233;
        test_data[2320] = 33'd2492348860;
        test_addr[2321] = 234;
        test_data[2321] = 33'd5638139681;
        test_addr[2322] = 235;
        test_data[2322] = 33'd597555204;
        test_addr[2323] = 236;
        test_data[2323] = 33'd2253456555;
        test_addr[2324] = 237;
        test_data[2324] = 33'd854297306;
        test_addr[2325] = 238;
        test_data[2325] = 33'd7377634913;
        test_addr[2326] = 239;
        test_data[2326] = 33'd6488619841;
        test_addr[2327] = 240;
        test_data[2327] = 33'd332704183;
        test_addr[2328] = 241;
        test_data[2328] = 33'd3112036660;
        test_addr[2329] = 242;
        test_data[2329] = 33'd7453344164;
        test_addr[2330] = 243;
        test_data[2330] = 33'd3483456815;
        test_addr[2331] = 87;
        test_data[2331] = 33'd1074381877;
        test_addr[2332] = 88;
        test_data[2332] = 33'd5149978986;
        test_addr[2333] = 89;
        test_data[2333] = 33'd3266191666;
        test_addr[2334] = 90;
        test_data[2334] = 33'd847785320;
        test_addr[2335] = 91;
        test_data[2335] = 33'd850272629;
        test_addr[2336] = 92;
        test_data[2336] = 33'd1952513095;
        test_addr[2337] = 93;
        test_data[2337] = 33'd2224978568;
        test_addr[2338] = 94;
        test_data[2338] = 33'd3836173812;
        test_addr[2339] = 95;
        test_data[2339] = 33'd3343865750;
        test_addr[2340] = 96;
        test_data[2340] = 33'd8326221411;
        test_addr[2341] = 97;
        test_data[2341] = 33'd5011617602;
        test_addr[2342] = 98;
        test_data[2342] = 33'd3796967958;
        test_addr[2343] = 99;
        test_data[2343] = 33'd3818727437;
        test_addr[2344] = 100;
        test_data[2344] = 33'd2034825318;
        test_addr[2345] = 101;
        test_data[2345] = 33'd352556074;
        test_addr[2346] = 102;
        test_data[2346] = 33'd736369780;
        test_addr[2347] = 103;
        test_data[2347] = 33'd7813199684;
        test_addr[2348] = 104;
        test_data[2348] = 33'd4549352016;
        test_addr[2349] = 105;
        test_data[2349] = 33'd3876404727;
        test_addr[2350] = 664;
        test_data[2350] = 33'd4123313617;
        test_addr[2351] = 665;
        test_data[2351] = 33'd8374910207;
        test_addr[2352] = 666;
        test_data[2352] = 33'd438118782;
        test_addr[2353] = 667;
        test_data[2353] = 33'd1504348005;
        test_addr[2354] = 668;
        test_data[2354] = 33'd7295078110;
        test_addr[2355] = 106;
        test_data[2355] = 33'd8102545914;
        test_addr[2356] = 107;
        test_data[2356] = 33'd3862762663;
        test_addr[2357] = 108;
        test_data[2357] = 33'd2831210998;
        test_addr[2358] = 109;
        test_data[2358] = 33'd7221713441;
        test_addr[2359] = 110;
        test_data[2359] = 33'd4423760897;
        test_addr[2360] = 111;
        test_data[2360] = 33'd6429036899;
        test_addr[2361] = 112;
        test_data[2361] = 33'd7690164071;
        test_addr[2362] = 113;
        test_data[2362] = 33'd958838625;
        test_addr[2363] = 114;
        test_data[2363] = 33'd2378794530;
        test_addr[2364] = 115;
        test_data[2364] = 33'd1652892941;
        test_addr[2365] = 116;
        test_data[2365] = 33'd2375022544;
        test_addr[2366] = 117;
        test_data[2366] = 33'd5950560693;
        test_addr[2367] = 118;
        test_data[2367] = 33'd6133224407;
        test_addr[2368] = 119;
        test_data[2368] = 33'd663222617;
        test_addr[2369] = 120;
        test_data[2369] = 33'd827454364;
        test_addr[2370] = 121;
        test_data[2370] = 33'd2605200182;
        test_addr[2371] = 122;
        test_data[2371] = 33'd3622924683;
        test_addr[2372] = 123;
        test_data[2372] = 33'd7747833304;
        test_addr[2373] = 35;
        test_data[2373] = 33'd1560223761;
        test_addr[2374] = 36;
        test_data[2374] = 33'd4012222965;
        test_addr[2375] = 37;
        test_data[2375] = 33'd2174070789;
        test_addr[2376] = 38;
        test_data[2376] = 33'd8459245881;
        test_addr[2377] = 39;
        test_data[2377] = 33'd407243807;
        test_addr[2378] = 40;
        test_data[2378] = 33'd5721084907;
        test_addr[2379] = 41;
        test_data[2379] = 33'd4778701022;
        test_addr[2380] = 42;
        test_data[2380] = 33'd6801386510;
        test_addr[2381] = 43;
        test_data[2381] = 33'd7078104309;
        test_addr[2382] = 124;
        test_data[2382] = 33'd7075738100;
        test_addr[2383] = 125;
        test_data[2383] = 33'd8089972385;
        test_addr[2384] = 126;
        test_data[2384] = 33'd989367641;
        test_addr[2385] = 127;
        test_data[2385] = 33'd972800406;
        test_addr[2386] = 128;
        test_data[2386] = 33'd8434026805;
        test_addr[2387] = 129;
        test_data[2387] = 33'd212359631;
        test_addr[2388] = 130;
        test_data[2388] = 33'd3185392084;
        test_addr[2389] = 925;
        test_data[2389] = 33'd3444626246;
        test_addr[2390] = 926;
        test_data[2390] = 33'd7353819508;
        test_addr[2391] = 927;
        test_data[2391] = 33'd4323355291;
        test_addr[2392] = 928;
        test_data[2392] = 33'd8526494587;
        test_addr[2393] = 131;
        test_data[2393] = 33'd2412978687;
        test_addr[2394] = 132;
        test_data[2394] = 33'd5192671196;
        test_addr[2395] = 133;
        test_data[2395] = 33'd1490977139;
        test_addr[2396] = 134;
        test_data[2396] = 33'd3657150815;
        test_addr[2397] = 135;
        test_data[2397] = 33'd7114671060;
        test_addr[2398] = 136;
        test_data[2398] = 33'd3351615148;
        test_addr[2399] = 137;
        test_data[2399] = 33'd3516062355;
        test_addr[2400] = 138;
        test_data[2400] = 33'd1254375529;
        test_addr[2401] = 866;
        test_data[2401] = 33'd636310232;
        test_addr[2402] = 867;
        test_data[2402] = 33'd4191967086;
        test_addr[2403] = 868;
        test_data[2403] = 33'd4926686794;
        test_addr[2404] = 869;
        test_data[2404] = 33'd6197803228;
        test_addr[2405] = 870;
        test_data[2405] = 33'd1319303959;
        test_addr[2406] = 871;
        test_data[2406] = 33'd7527389338;
        test_addr[2407] = 872;
        test_data[2407] = 33'd3833194746;
        test_addr[2408] = 139;
        test_data[2408] = 33'd4040208455;
        test_addr[2409] = 140;
        test_data[2409] = 33'd452007419;
        test_addr[2410] = 141;
        test_data[2410] = 33'd7981335879;
        test_addr[2411] = 142;
        test_data[2411] = 33'd2878388451;
        test_addr[2412] = 143;
        test_data[2412] = 33'd7715034;
        test_addr[2413] = 144;
        test_data[2413] = 33'd1365519167;
        test_addr[2414] = 145;
        test_data[2414] = 33'd2955818252;
        test_addr[2415] = 564;
        test_data[2415] = 33'd869541130;
        test_addr[2416] = 565;
        test_data[2416] = 33'd1714782340;
        test_addr[2417] = 566;
        test_data[2417] = 33'd2303519254;
        test_addr[2418] = 146;
        test_data[2418] = 33'd111211454;
        test_addr[2419] = 147;
        test_data[2419] = 33'd8583594589;
        test_addr[2420] = 148;
        test_data[2420] = 33'd6952297730;
        test_addr[2421] = 149;
        test_data[2421] = 33'd5171649377;
        test_addr[2422] = 150;
        test_data[2422] = 33'd1569648152;
        test_addr[2423] = 151;
        test_data[2423] = 33'd1553933429;
        test_addr[2424] = 152;
        test_data[2424] = 33'd2253932096;
        test_addr[2425] = 153;
        test_data[2425] = 33'd3061874645;
        test_addr[2426] = 154;
        test_data[2426] = 33'd8184554214;
        test_addr[2427] = 155;
        test_data[2427] = 33'd8029931863;
        test_addr[2428] = 156;
        test_data[2428] = 33'd6956058983;
        test_addr[2429] = 157;
        test_data[2429] = 33'd2310668724;
        test_addr[2430] = 158;
        test_data[2430] = 33'd3556418516;
        test_addr[2431] = 159;
        test_data[2431] = 33'd3037698070;
        test_addr[2432] = 160;
        test_data[2432] = 33'd7697581497;
        test_addr[2433] = 161;
        test_data[2433] = 33'd4580329586;
        test_addr[2434] = 162;
        test_data[2434] = 33'd3143417896;
        test_addr[2435] = 163;
        test_data[2435] = 33'd3528470030;
        test_addr[2436] = 164;
        test_data[2436] = 33'd342696692;
        test_addr[2437] = 672;
        test_data[2437] = 33'd7644459037;
        test_addr[2438] = 673;
        test_data[2438] = 33'd7264629088;
        test_addr[2439] = 674;
        test_data[2439] = 33'd1684633886;
        test_addr[2440] = 675;
        test_data[2440] = 33'd3494862483;
        test_addr[2441] = 676;
        test_data[2441] = 33'd662578081;
        test_addr[2442] = 677;
        test_data[2442] = 33'd1877633440;
        test_addr[2443] = 678;
        test_data[2443] = 33'd4202950769;
        test_addr[2444] = 679;
        test_data[2444] = 33'd2237167224;
        test_addr[2445] = 680;
        test_data[2445] = 33'd8504883541;
        test_addr[2446] = 681;
        test_data[2446] = 33'd3197818006;
        test_addr[2447] = 682;
        test_data[2447] = 33'd666405120;
        test_addr[2448] = 683;
        test_data[2448] = 33'd1731237928;
        test_addr[2449] = 165;
        test_data[2449] = 33'd3597588474;
        test_addr[2450] = 166;
        test_data[2450] = 33'd2253906058;
        test_addr[2451] = 167;
        test_data[2451] = 33'd367704174;
        test_addr[2452] = 168;
        test_data[2452] = 33'd864052885;
        test_addr[2453] = 169;
        test_data[2453] = 33'd3020898125;
        test_addr[2454] = 91;
        test_data[2454] = 33'd850272629;
        test_addr[2455] = 92;
        test_data[2455] = 33'd1952513095;
        test_addr[2456] = 93;
        test_data[2456] = 33'd2224978568;
        test_addr[2457] = 94;
        test_data[2457] = 33'd3836173812;
        test_addr[2458] = 95;
        test_data[2458] = 33'd5248806697;
        test_addr[2459] = 96;
        test_data[2459] = 33'd4031254115;
        test_addr[2460] = 97;
        test_data[2460] = 33'd716650306;
        test_addr[2461] = 98;
        test_data[2461] = 33'd3796967958;
        test_addr[2462] = 99;
        test_data[2462] = 33'd3818727437;
        test_addr[2463] = 100;
        test_data[2463] = 33'd2034825318;
        test_addr[2464] = 101;
        test_data[2464] = 33'd352556074;
        test_addr[2465] = 102;
        test_data[2465] = 33'd7573606898;
        test_addr[2466] = 103;
        test_data[2466] = 33'd3518232388;
        test_addr[2467] = 104;
        test_data[2467] = 33'd254384720;
        test_addr[2468] = 105;
        test_data[2468] = 33'd3876404727;
        test_addr[2469] = 106;
        test_data[2469] = 33'd3807578618;
        test_addr[2470] = 107;
        test_data[2470] = 33'd3862762663;
        test_addr[2471] = 108;
        test_data[2471] = 33'd4811642516;
        test_addr[2472] = 109;
        test_data[2472] = 33'd2926746145;
        test_addr[2473] = 170;
        test_data[2473] = 33'd911045719;
        test_addr[2474] = 171;
        test_data[2474] = 33'd4210643370;
        test_addr[2475] = 172;
        test_data[2475] = 33'd3645680872;
        test_addr[2476] = 173;
        test_data[2476] = 33'd7756667019;
        test_addr[2477] = 844;
        test_data[2477] = 33'd7924544170;
        test_addr[2478] = 845;
        test_data[2478] = 33'd6584526485;
        test_addr[2479] = 846;
        test_data[2479] = 33'd3129315442;
        test_addr[2480] = 847;
        test_data[2480] = 33'd5815542621;
        test_addr[2481] = 848;
        test_data[2481] = 33'd8379565311;
        test_addr[2482] = 849;
        test_data[2482] = 33'd4088205861;
        test_addr[2483] = 850;
        test_data[2483] = 33'd3650411410;
        test_addr[2484] = 851;
        test_data[2484] = 33'd8191170286;
        test_addr[2485] = 852;
        test_data[2485] = 33'd2704192971;
        test_addr[2486] = 853;
        test_data[2486] = 33'd1067052146;
        test_addr[2487] = 854;
        test_data[2487] = 33'd7096307341;
        test_addr[2488] = 855;
        test_data[2488] = 33'd5899502141;
        test_addr[2489] = 174;
        test_data[2489] = 33'd1152654674;
        test_addr[2490] = 175;
        test_data[2490] = 33'd5551226381;
        test_addr[2491] = 484;
        test_data[2491] = 33'd998179708;
        test_addr[2492] = 485;
        test_data[2492] = 33'd1497784997;
        test_addr[2493] = 486;
        test_data[2493] = 33'd7150131889;
        test_addr[2494] = 487;
        test_data[2494] = 33'd4233924408;
        test_addr[2495] = 488;
        test_data[2495] = 33'd3230286556;
        test_addr[2496] = 489;
        test_data[2496] = 33'd7602361293;
        test_addr[2497] = 176;
        test_data[2497] = 33'd3906597641;
        test_addr[2498] = 177;
        test_data[2498] = 33'd8405311329;
        test_addr[2499] = 178;
        test_data[2499] = 33'd3878152893;
        test_addr[2500] = 179;
        test_data[2500] = 33'd4900149937;
        test_addr[2501] = 180;
        test_data[2501] = 33'd5280967633;
        test_addr[2502] = 181;
        test_data[2502] = 33'd4739030047;
        test_addr[2503] = 182;
        test_data[2503] = 33'd3172527317;
        test_addr[2504] = 183;
        test_data[2504] = 33'd792941705;
        test_addr[2505] = 184;
        test_data[2505] = 33'd6223845061;
        test_addr[2506] = 185;
        test_data[2506] = 33'd2391399405;
        test_addr[2507] = 186;
        test_data[2507] = 33'd3062031139;
        test_addr[2508] = 187;
        test_data[2508] = 33'd793217816;
        test_addr[2509] = 188;
        test_data[2509] = 33'd8580644526;
        test_addr[2510] = 189;
        test_data[2510] = 33'd2741390496;
        test_addr[2511] = 190;
        test_data[2511] = 33'd3674547407;
        test_addr[2512] = 501;
        test_data[2512] = 33'd2592532499;
        test_addr[2513] = 502;
        test_data[2513] = 33'd1661402023;
        test_addr[2514] = 503;
        test_data[2514] = 33'd1739400798;
        test_addr[2515] = 504;
        test_data[2515] = 33'd225331988;
        test_addr[2516] = 505;
        test_data[2516] = 33'd977986578;
        test_addr[2517] = 506;
        test_data[2517] = 33'd7604852669;
        test_addr[2518] = 507;
        test_data[2518] = 33'd3984605869;
        test_addr[2519] = 508;
        test_data[2519] = 33'd1247575968;
        test_addr[2520] = 191;
        test_data[2520] = 33'd7340244519;
        test_addr[2521] = 192;
        test_data[2521] = 33'd5072378689;
        test_addr[2522] = 193;
        test_data[2522] = 33'd1033777528;
        test_addr[2523] = 194;
        test_data[2523] = 33'd2955644450;
        test_addr[2524] = 195;
        test_data[2524] = 33'd2193846095;
        test_addr[2525] = 196;
        test_data[2525] = 33'd2584950764;
        test_addr[2526] = 197;
        test_data[2526] = 33'd1696743885;
        test_addr[2527] = 198;
        test_data[2527] = 33'd2875093575;
        test_addr[2528] = 199;
        test_data[2528] = 33'd117868309;
        test_addr[2529] = 200;
        test_data[2529] = 33'd4066794897;
        test_addr[2530] = 201;
        test_data[2530] = 33'd1479348861;
        test_addr[2531] = 202;
        test_data[2531] = 33'd6186435425;
        test_addr[2532] = 203;
        test_data[2532] = 33'd8386683781;
        test_addr[2533] = 204;
        test_data[2533] = 33'd4344654462;
        test_addr[2534] = 205;
        test_data[2534] = 33'd382451800;
        test_addr[2535] = 206;
        test_data[2535] = 33'd4213338333;
        test_addr[2536] = 207;
        test_data[2536] = 33'd513445133;
        test_addr[2537] = 208;
        test_data[2537] = 33'd6374911225;
        test_addr[2538] = 209;
        test_data[2538] = 33'd3259078447;
        test_addr[2539] = 210;
        test_data[2539] = 33'd118596569;
        test_addr[2540] = 244;
        test_data[2540] = 33'd7074652529;
        test_addr[2541] = 245;
        test_data[2541] = 33'd4596019133;
        test_addr[2542] = 246;
        test_data[2542] = 33'd5138885097;
        test_addr[2543] = 247;
        test_data[2543] = 33'd3793934249;
        test_addr[2544] = 248;
        test_data[2544] = 33'd908055748;
        test_addr[2545] = 249;
        test_data[2545] = 33'd3317083412;
        test_addr[2546] = 250;
        test_data[2546] = 33'd6910404597;
        test_addr[2547] = 251;
        test_data[2547] = 33'd5782342842;
        test_addr[2548] = 252;
        test_data[2548] = 33'd855026393;
        test_addr[2549] = 253;
        test_data[2549] = 33'd2844318793;
        test_addr[2550] = 211;
        test_data[2550] = 33'd4202191155;
        test_addr[2551] = 315;
        test_data[2551] = 33'd7091404319;
        test_addr[2552] = 316;
        test_data[2552] = 33'd4113165209;
        test_addr[2553] = 317;
        test_data[2553] = 33'd2374556068;
        test_addr[2554] = 318;
        test_data[2554] = 33'd1665876031;
        test_addr[2555] = 319;
        test_data[2555] = 33'd5953829139;
        test_addr[2556] = 212;
        test_data[2556] = 33'd2809482033;
        test_addr[2557] = 1;
        test_data[2557] = 33'd6164542229;
        test_addr[2558] = 2;
        test_data[2558] = 33'd728813621;
        test_addr[2559] = 3;
        test_data[2559] = 33'd2095642455;
        test_addr[2560] = 4;
        test_data[2560] = 33'd925613716;
        test_addr[2561] = 5;
        test_data[2561] = 33'd485978242;
        test_addr[2562] = 6;
        test_data[2562] = 33'd5449070952;
        test_addr[2563] = 7;
        test_data[2563] = 33'd966600747;
        test_addr[2564] = 8;
        test_data[2564] = 33'd3378399337;
        test_addr[2565] = 9;
        test_data[2565] = 33'd5409008510;
        test_addr[2566] = 10;
        test_data[2566] = 33'd7844920347;
        test_addr[2567] = 11;
        test_data[2567] = 33'd5169814738;
        test_addr[2568] = 12;
        test_data[2568] = 33'd1442523325;
        test_addr[2569] = 213;
        test_data[2569] = 33'd3848169259;
        test_addr[2570] = 214;
        test_data[2570] = 33'd635033231;
        test_addr[2571] = 215;
        test_data[2571] = 33'd4098659685;
        test_addr[2572] = 216;
        test_data[2572] = 33'd1581642574;
        test_addr[2573] = 217;
        test_data[2573] = 33'd2718828492;
        test_addr[2574] = 218;
        test_data[2574] = 33'd7568580299;
        test_addr[2575] = 219;
        test_data[2575] = 33'd1518323074;
        test_addr[2576] = 220;
        test_data[2576] = 33'd5307350323;
        test_addr[2577] = 221;
        test_data[2577] = 33'd3019464660;
        test_addr[2578] = 146;
        test_data[2578] = 33'd7468799338;
        test_addr[2579] = 147;
        test_data[2579] = 33'd4288627293;
        test_addr[2580] = 148;
        test_data[2580] = 33'd5387855751;
        test_addr[2581] = 149;
        test_data[2581] = 33'd876682081;
        test_addr[2582] = 150;
        test_data[2582] = 33'd6753423962;
        test_addr[2583] = 151;
        test_data[2583] = 33'd1553933429;
        test_addr[2584] = 152;
        test_data[2584] = 33'd2253932096;
        test_addr[2585] = 153;
        test_data[2585] = 33'd3061874645;
        test_addr[2586] = 154;
        test_data[2586] = 33'd7550049105;
        test_addr[2587] = 155;
        test_data[2587] = 33'd5163594214;
        test_addr[2588] = 222;
        test_data[2588] = 33'd1384897455;
        test_addr[2589] = 223;
        test_data[2589] = 33'd5564601043;
        test_addr[2590] = 224;
        test_data[2590] = 33'd4539215933;
        test_addr[2591] = 225;
        test_data[2591] = 33'd1457651049;
        test_addr[2592] = 226;
        test_data[2592] = 33'd3315378073;
        test_addr[2593] = 227;
        test_data[2593] = 33'd2688484918;
        test_addr[2594] = 228;
        test_data[2594] = 33'd4120475529;
        test_addr[2595] = 229;
        test_data[2595] = 33'd5454082161;
        test_addr[2596] = 230;
        test_data[2596] = 33'd988458485;
        test_addr[2597] = 231;
        test_data[2597] = 33'd6551801561;
        test_addr[2598] = 232;
        test_data[2598] = 33'd5377065558;
        test_addr[2599] = 90;
        test_data[2599] = 33'd5519377413;
        test_addr[2600] = 91;
        test_data[2600] = 33'd850272629;
        test_addr[2601] = 92;
        test_data[2601] = 33'd1952513095;
        test_addr[2602] = 93;
        test_data[2602] = 33'd2224978568;
        test_addr[2603] = 94;
        test_data[2603] = 33'd7574141903;
        test_addr[2604] = 95;
        test_data[2604] = 33'd953839401;
        test_addr[2605] = 96;
        test_data[2605] = 33'd4031254115;
        test_addr[2606] = 97;
        test_data[2606] = 33'd8468470577;
        test_addr[2607] = 98;
        test_data[2607] = 33'd4980207096;
        test_addr[2608] = 99;
        test_data[2608] = 33'd6179235705;
        test_addr[2609] = 100;
        test_data[2609] = 33'd6374626038;
        test_addr[2610] = 101;
        test_data[2610] = 33'd6028492966;
        test_addr[2611] = 233;
        test_data[2611] = 33'd5933643083;
        test_addr[2612] = 234;
        test_data[2612] = 33'd4746574840;
        test_addr[2613] = 235;
        test_data[2613] = 33'd597555204;
        test_addr[2614] = 236;
        test_data[2614] = 33'd7393604384;
        test_addr[2615] = 237;
        test_data[2615] = 33'd854297306;
        test_addr[2616] = 238;
        test_data[2616] = 33'd3082667617;
        test_addr[2617] = 239;
        test_data[2617] = 33'd6173207494;
        test_addr[2618] = 240;
        test_data[2618] = 33'd332704183;
        test_addr[2619] = 359;
        test_data[2619] = 33'd3907129635;
        test_addr[2620] = 360;
        test_data[2620] = 33'd202881912;
        test_addr[2621] = 361;
        test_data[2621] = 33'd2414551097;
        test_addr[2622] = 362;
        test_data[2622] = 33'd7963468466;
        test_addr[2623] = 363;
        test_data[2623] = 33'd2723076636;
        test_addr[2624] = 364;
        test_data[2624] = 33'd1333182938;
        test_addr[2625] = 365;
        test_data[2625] = 33'd1161783265;
        test_addr[2626] = 366;
        test_data[2626] = 33'd7208775220;
        test_addr[2627] = 367;
        test_data[2627] = 33'd3426483264;
        test_addr[2628] = 368;
        test_data[2628] = 33'd384401585;
        test_addr[2629] = 369;
        test_data[2629] = 33'd2107994983;
        test_addr[2630] = 241;
        test_data[2630] = 33'd3112036660;
        test_addr[2631] = 242;
        test_data[2631] = 33'd5215431782;
        test_addr[2632] = 243;
        test_data[2632] = 33'd3483456815;
        test_addr[2633] = 244;
        test_data[2633] = 33'd2779685233;
        test_addr[2634] = 245;
        test_data[2634] = 33'd301051837;
        test_addr[2635] = 246;
        test_data[2635] = 33'd6185684529;
        test_addr[2636] = 247;
        test_data[2636] = 33'd3793934249;
        test_addr[2637] = 248;
        test_data[2637] = 33'd908055748;
        test_addr[2638] = 249;
        test_data[2638] = 33'd7486029019;
        test_addr[2639] = 250;
        test_data[2639] = 33'd2615437301;
        test_addr[2640] = 251;
        test_data[2640] = 33'd1487375546;
        test_addr[2641] = 252;
        test_data[2641] = 33'd4539018454;
        test_addr[2642] = 253;
        test_data[2642] = 33'd8518729367;
        test_addr[2643] = 254;
        test_data[2643] = 33'd100893370;
        test_addr[2644] = 255;
        test_data[2644] = 33'd2507835843;
        test_addr[2645] = 256;
        test_data[2645] = 33'd4960430147;
        test_addr[2646] = 257;
        test_data[2646] = 33'd4311298278;
        test_addr[2647] = 258;
        test_data[2647] = 33'd1463838338;
        test_addr[2648] = 259;
        test_data[2648] = 33'd5422308072;
        test_addr[2649] = 260;
        test_data[2649] = 33'd7104130718;
        test_addr[2650] = 261;
        test_data[2650] = 33'd4986471997;
        test_addr[2651] = 224;
        test_data[2651] = 33'd244248637;
        test_addr[2652] = 225;
        test_data[2652] = 33'd6900608531;
        test_addr[2653] = 226;
        test_data[2653] = 33'd5861400700;
        test_addr[2654] = 227;
        test_data[2654] = 33'd2688484918;
        test_addr[2655] = 228;
        test_data[2655] = 33'd8339031550;
        test_addr[2656] = 229;
        test_data[2656] = 33'd1159114865;
        test_addr[2657] = 262;
        test_data[2657] = 33'd3224676958;
        test_addr[2658] = 263;
        test_data[2658] = 33'd3200855956;
        test_addr[2659] = 264;
        test_data[2659] = 33'd4124826968;
        test_addr[2660] = 265;
        test_data[2660] = 33'd2848828629;
        test_addr[2661] = 266;
        test_data[2661] = 33'd2745001205;
        test_addr[2662] = 267;
        test_data[2662] = 33'd5388337768;
        test_addr[2663] = 268;
        test_data[2663] = 33'd189083836;
        test_addr[2664] = 269;
        test_data[2664] = 33'd90054363;
        test_addr[2665] = 270;
        test_data[2665] = 33'd4155868294;
        test_addr[2666] = 271;
        test_data[2666] = 33'd6303686877;
        test_addr[2667] = 272;
        test_data[2667] = 33'd7560741678;
        test_addr[2668] = 273;
        test_data[2668] = 33'd5398244738;
        test_addr[2669] = 274;
        test_data[2669] = 33'd5895128397;
        test_addr[2670] = 275;
        test_data[2670] = 33'd1254626076;
        test_addr[2671] = 498;
        test_data[2671] = 33'd4163492510;
        test_addr[2672] = 499;
        test_data[2672] = 33'd5126442863;
        test_addr[2673] = 276;
        test_data[2673] = 33'd2468941697;
        test_addr[2674] = 277;
        test_data[2674] = 33'd1644482855;
        test_addr[2675] = 278;
        test_data[2675] = 33'd1532905441;
        test_addr[2676] = 279;
        test_data[2676] = 33'd4221166951;
        test_addr[2677] = 280;
        test_data[2677] = 33'd924432628;
        test_addr[2678] = 281;
        test_data[2678] = 33'd6826022249;
        test_addr[2679] = 282;
        test_data[2679] = 33'd7938480391;
        test_addr[2680] = 283;
        test_data[2680] = 33'd7833730974;
        test_addr[2681] = 284;
        test_data[2681] = 33'd5459348886;
        test_addr[2682] = 285;
        test_data[2682] = 33'd3139190243;
        test_addr[2683] = 286;
        test_data[2683] = 33'd2132904872;
        test_addr[2684] = 287;
        test_data[2684] = 33'd4288613521;
        test_addr[2685] = 288;
        test_data[2685] = 33'd6824259681;
        test_addr[2686] = 289;
        test_data[2686] = 33'd7392686736;
        test_addr[2687] = 290;
        test_data[2687] = 33'd2038912635;
        test_addr[2688] = 291;
        test_data[2688] = 33'd2507289981;
        test_addr[2689] = 292;
        test_data[2689] = 33'd1640016259;
        test_addr[2690] = 293;
        test_data[2690] = 33'd1249044169;
        test_addr[2691] = 294;
        test_data[2691] = 33'd7363543031;
        test_addr[2692] = 295;
        test_data[2692] = 33'd6721086909;
        test_addr[2693] = 296;
        test_data[2693] = 33'd366076987;
        test_addr[2694] = 297;
        test_data[2694] = 33'd2331663310;
        test_addr[2695] = 298;
        test_data[2695] = 33'd724689699;
        test_addr[2696] = 299;
        test_data[2696] = 33'd5909302975;
        test_addr[2697] = 300;
        test_data[2697] = 33'd5357910562;
        test_addr[2698] = 603;
        test_data[2698] = 33'd2792617507;
        test_addr[2699] = 604;
        test_data[2699] = 33'd998324771;
        test_addr[2700] = 605;
        test_data[2700] = 33'd1618144234;
        test_addr[2701] = 606;
        test_data[2701] = 33'd920782161;
        test_addr[2702] = 607;
        test_data[2702] = 33'd3986635328;
        test_addr[2703] = 608;
        test_data[2703] = 33'd2953791377;
        test_addr[2704] = 609;
        test_data[2704] = 33'd6869915917;
        test_addr[2705] = 610;
        test_data[2705] = 33'd4895450635;
        test_addr[2706] = 611;
        test_data[2706] = 33'd6359124314;
        test_addr[2707] = 612;
        test_data[2707] = 33'd3706301070;
        test_addr[2708] = 613;
        test_data[2708] = 33'd1070746388;
        test_addr[2709] = 614;
        test_data[2709] = 33'd2106134210;
        test_addr[2710] = 615;
        test_data[2710] = 33'd7131505305;
        test_addr[2711] = 616;
        test_data[2711] = 33'd2279850305;
        test_addr[2712] = 301;
        test_data[2712] = 33'd3116504789;
        test_addr[2713] = 302;
        test_data[2713] = 33'd3657246985;
        test_addr[2714] = 214;
        test_data[2714] = 33'd8518369902;
        test_addr[2715] = 215;
        test_data[2715] = 33'd4098659685;
        test_addr[2716] = 216;
        test_data[2716] = 33'd1581642574;
        test_addr[2717] = 217;
        test_data[2717] = 33'd2718828492;
        test_addr[2718] = 218;
        test_data[2718] = 33'd3273613003;
        test_addr[2719] = 219;
        test_data[2719] = 33'd1518323074;
        test_addr[2720] = 220;
        test_data[2720] = 33'd1012383027;
        test_addr[2721] = 221;
        test_data[2721] = 33'd3019464660;
        test_addr[2722] = 222;
        test_data[2722] = 33'd1384897455;
        test_addr[2723] = 223;
        test_data[2723] = 33'd5883857258;
        test_addr[2724] = 224;
        test_data[2724] = 33'd6426310932;
        test_addr[2725] = 225;
        test_data[2725] = 33'd2605641235;
        test_addr[2726] = 226;
        test_data[2726] = 33'd5721209928;
        test_addr[2727] = 227;
        test_data[2727] = 33'd5030493555;
        test_addr[2728] = 228;
        test_data[2728] = 33'd4044064254;
        test_addr[2729] = 229;
        test_data[2729] = 33'd1159114865;
        test_addr[2730] = 230;
        test_data[2730] = 33'd988458485;
        test_addr[2731] = 231;
        test_data[2731] = 33'd2256834265;
        test_addr[2732] = 232;
        test_data[2732] = 33'd1082098262;
        test_addr[2733] = 303;
        test_data[2733] = 33'd6434928683;
        test_addr[2734] = 304;
        test_data[2734] = 33'd3620887989;
        test_addr[2735] = 305;
        test_data[2735] = 33'd3296594168;
        test_addr[2736] = 306;
        test_data[2736] = 33'd3900608396;
        test_addr[2737] = 307;
        test_data[2737] = 33'd144487780;
        test_addr[2738] = 935;
        test_data[2738] = 33'd2918620527;
        test_addr[2739] = 936;
        test_data[2739] = 33'd7932397066;
        test_addr[2740] = 937;
        test_data[2740] = 33'd1191377286;
        test_addr[2741] = 938;
        test_data[2741] = 33'd5096224200;
        test_addr[2742] = 939;
        test_data[2742] = 33'd775116840;
        test_addr[2743] = 940;
        test_data[2743] = 33'd3766189908;
        test_addr[2744] = 941;
        test_data[2744] = 33'd4232471274;
        test_addr[2745] = 942;
        test_data[2745] = 33'd7576008826;
        test_addr[2746] = 943;
        test_data[2746] = 33'd7479496002;
        test_addr[2747] = 308;
        test_data[2747] = 33'd315191869;
        test_addr[2748] = 123;
        test_data[2748] = 33'd3452866008;
        test_addr[2749] = 309;
        test_data[2749] = 33'd7079933450;
        test_addr[2750] = 310;
        test_data[2750] = 33'd727353973;
        test_addr[2751] = 311;
        test_data[2751] = 33'd4814452369;
        test_addr[2752] = 312;
        test_data[2752] = 33'd6488838379;
        test_addr[2753] = 313;
        test_data[2753] = 33'd2458964169;
        test_addr[2754] = 314;
        test_data[2754] = 33'd8286379279;
        test_addr[2755] = 315;
        test_data[2755] = 33'd5708679611;
        test_addr[2756] = 316;
        test_data[2756] = 33'd4113165209;
        test_addr[2757] = 82;
        test_data[2757] = 33'd6074193997;
        test_addr[2758] = 317;
        test_data[2758] = 33'd2374556068;
        test_addr[2759] = 318;
        test_data[2759] = 33'd1665876031;
        test_addr[2760] = 114;
        test_data[2760] = 33'd2378794530;
        test_addr[2761] = 115;
        test_data[2761] = 33'd4362308329;
        test_addr[2762] = 116;
        test_data[2762] = 33'd2375022544;
        test_addr[2763] = 117;
        test_data[2763] = 33'd1655593397;
        test_addr[2764] = 118;
        test_data[2764] = 33'd5424234904;
        test_addr[2765] = 119;
        test_data[2765] = 33'd663222617;
        test_addr[2766] = 120;
        test_data[2766] = 33'd827454364;
        test_addr[2767] = 121;
        test_data[2767] = 33'd2605200182;
        test_addr[2768] = 122;
        test_data[2768] = 33'd3622924683;
        test_addr[2769] = 123;
        test_data[2769] = 33'd3452866008;
        test_addr[2770] = 124;
        test_data[2770] = 33'd2780770804;
        test_addr[2771] = 125;
        test_data[2771] = 33'd4347929018;
        test_addr[2772] = 126;
        test_data[2772] = 33'd8485429833;
        test_addr[2773] = 127;
        test_data[2773] = 33'd972800406;
        test_addr[2774] = 128;
        test_data[2774] = 33'd4139059509;
        test_addr[2775] = 129;
        test_data[2775] = 33'd212359631;
        test_addr[2776] = 130;
        test_data[2776] = 33'd4667438569;
        test_addr[2777] = 131;
        test_data[2777] = 33'd2412978687;
        test_addr[2778] = 132;
        test_data[2778] = 33'd6577082798;
        test_addr[2779] = 133;
        test_data[2779] = 33'd1490977139;
        test_addr[2780] = 134;
        test_data[2780] = 33'd3657150815;
        test_addr[2781] = 135;
        test_data[2781] = 33'd2819703764;
        test_addr[2782] = 136;
        test_data[2782] = 33'd3351615148;
        test_addr[2783] = 137;
        test_data[2783] = 33'd3516062355;
        test_addr[2784] = 138;
        test_data[2784] = 33'd1254375529;
        test_addr[2785] = 139;
        test_data[2785] = 33'd7593361222;
        test_addr[2786] = 319;
        test_data[2786] = 33'd6515735976;
        test_addr[2787] = 916;
        test_data[2787] = 33'd5212806837;
        test_addr[2788] = 917;
        test_data[2788] = 33'd7878205887;
        test_addr[2789] = 918;
        test_data[2789] = 33'd771796738;
        test_addr[2790] = 320;
        test_data[2790] = 33'd2364460379;
        test_addr[2791] = 321;
        test_data[2791] = 33'd4278979725;
        test_addr[2792] = 322;
        test_data[2792] = 33'd341336502;
        test_addr[2793] = 323;
        test_data[2793] = 33'd1953799233;
        test_addr[2794] = 324;
        test_data[2794] = 33'd8096359894;
        test_addr[2795] = 325;
        test_data[2795] = 33'd6480144236;
        test_addr[2796] = 326;
        test_data[2796] = 33'd586463684;
        test_addr[2797] = 327;
        test_data[2797] = 33'd739327056;
        test_addr[2798] = 328;
        test_data[2798] = 33'd2908366129;
        test_addr[2799] = 329;
        test_data[2799] = 33'd2309989022;
        test_addr[2800] = 330;
        test_data[2800] = 33'd3508612389;
        test_addr[2801] = 331;
        test_data[2801] = 33'd4229591735;
        test_addr[2802] = 332;
        test_data[2802] = 33'd4266769130;
        test_addr[2803] = 333;
        test_data[2803] = 33'd2296982685;
        test_addr[2804] = 334;
        test_data[2804] = 33'd1942623992;
        test_addr[2805] = 335;
        test_data[2805] = 33'd1195626943;
        test_addr[2806] = 336;
        test_data[2806] = 33'd1688024943;
        test_addr[2807] = 851;
        test_data[2807] = 33'd3896202990;
        test_addr[2808] = 852;
        test_data[2808] = 33'd2704192971;
        test_addr[2809] = 853;
        test_data[2809] = 33'd1067052146;
        test_addr[2810] = 337;
        test_data[2810] = 33'd750261429;
        test_addr[2811] = 338;
        test_data[2811] = 33'd1821314294;
        test_addr[2812] = 339;
        test_data[2812] = 33'd3966375939;
        test_addr[2813] = 340;
        test_data[2813] = 33'd5683974501;
        test_addr[2814] = 341;
        test_data[2814] = 33'd315843574;
        test_addr[2815] = 342;
        test_data[2815] = 33'd421435128;
        test_addr[2816] = 343;
        test_data[2816] = 33'd2846218665;
        test_addr[2817] = 344;
        test_data[2817] = 33'd768223443;
        test_addr[2818] = 345;
        test_data[2818] = 33'd2791959723;
        test_addr[2819] = 346;
        test_data[2819] = 33'd6271636085;
        test_addr[2820] = 347;
        test_data[2820] = 33'd4150740891;
        test_addr[2821] = 348;
        test_data[2821] = 33'd7215780248;
        test_addr[2822] = 349;
        test_data[2822] = 33'd8416215247;
        test_addr[2823] = 350;
        test_data[2823] = 33'd6762763702;
        test_addr[2824] = 351;
        test_data[2824] = 33'd705076357;
        test_addr[2825] = 352;
        test_data[2825] = 33'd4515401125;
        test_addr[2826] = 353;
        test_data[2826] = 33'd2990531551;
        test_addr[2827] = 354;
        test_data[2827] = 33'd4080977870;
        test_addr[2828] = 355;
        test_data[2828] = 33'd2975558951;
        test_addr[2829] = 356;
        test_data[2829] = 33'd2257235136;
        test_addr[2830] = 357;
        test_data[2830] = 33'd4115832282;
        test_addr[2831] = 34;
        test_data[2831] = 33'd1469107037;
        test_addr[2832] = 35;
        test_data[2832] = 33'd1560223761;
        test_addr[2833] = 36;
        test_data[2833] = 33'd7620757408;
        test_addr[2834] = 358;
        test_data[2834] = 33'd5196125499;
        test_addr[2835] = 359;
        test_data[2835] = 33'd3907129635;
        test_addr[2836] = 360;
        test_data[2836] = 33'd202881912;
        test_addr[2837] = 361;
        test_data[2837] = 33'd2414551097;
        test_addr[2838] = 362;
        test_data[2838] = 33'd8279690572;
        test_addr[2839] = 363;
        test_data[2839] = 33'd2723076636;
        test_addr[2840] = 364;
        test_data[2840] = 33'd6009097462;
        test_addr[2841] = 534;
        test_data[2841] = 33'd2666228914;
        test_addr[2842] = 535;
        test_data[2842] = 33'd5920267521;
        test_addr[2843] = 536;
        test_data[2843] = 33'd979101880;
        test_addr[2844] = 537;
        test_data[2844] = 33'd1269482248;
        test_addr[2845] = 538;
        test_data[2845] = 33'd5470758519;
        test_addr[2846] = 539;
        test_data[2846] = 33'd1252831804;
        test_addr[2847] = 540;
        test_data[2847] = 33'd3769408227;
        test_addr[2848] = 541;
        test_data[2848] = 33'd6343915741;
        test_addr[2849] = 542;
        test_data[2849] = 33'd1354020355;
        test_addr[2850] = 543;
        test_data[2850] = 33'd4695240909;
        test_addr[2851] = 544;
        test_data[2851] = 33'd2499634813;
        test_addr[2852] = 545;
        test_data[2852] = 33'd8149817109;
        test_addr[2853] = 546;
        test_data[2853] = 33'd3953366411;
        test_addr[2854] = 547;
        test_data[2854] = 33'd2783941199;
        test_addr[2855] = 548;
        test_data[2855] = 33'd4827155212;
        test_addr[2856] = 549;
        test_data[2856] = 33'd2114883172;
        test_addr[2857] = 550;
        test_data[2857] = 33'd5361410940;
        test_addr[2858] = 551;
        test_data[2858] = 33'd3755615061;
        test_addr[2859] = 365;
        test_data[2859] = 33'd1161783265;
        test_addr[2860] = 366;
        test_data[2860] = 33'd5884553772;
        test_addr[2861] = 367;
        test_data[2861] = 33'd3426483264;
        test_addr[2862] = 552;
        test_data[2862] = 33'd2229852656;
        test_addr[2863] = 553;
        test_data[2863] = 33'd3462769718;
        test_addr[2864] = 554;
        test_data[2864] = 33'd717641719;
        test_addr[2865] = 555;
        test_data[2865] = 33'd3459416445;
        test_addr[2866] = 556;
        test_data[2866] = 33'd7164712655;
        test_addr[2867] = 557;
        test_data[2867] = 33'd5735740813;
        test_addr[2868] = 558;
        test_data[2868] = 33'd1593008829;
        test_addr[2869] = 559;
        test_data[2869] = 33'd1691044550;
        test_addr[2870] = 368;
        test_data[2870] = 33'd7449180479;
        test_addr[2871] = 369;
        test_data[2871] = 33'd2107994983;
        test_addr[2872] = 370;
        test_data[2872] = 33'd151832112;
        test_addr[2873] = 371;
        test_data[2873] = 33'd2775974076;
        test_addr[2874] = 372;
        test_data[2874] = 33'd6775323877;
        test_addr[2875] = 373;
        test_data[2875] = 33'd6443286441;
        test_addr[2876] = 374;
        test_data[2876] = 33'd4082071206;
        test_addr[2877] = 375;
        test_data[2877] = 33'd2719622023;
        test_addr[2878] = 376;
        test_data[2878] = 33'd7709473257;
        test_addr[2879] = 377;
        test_data[2879] = 33'd436835430;
        test_addr[2880] = 378;
        test_data[2880] = 33'd7915869209;
        test_addr[2881] = 379;
        test_data[2881] = 33'd708784957;
        test_addr[2882] = 380;
        test_data[2882] = 33'd5909915487;
        test_addr[2883] = 381;
        test_data[2883] = 33'd1741094807;
        test_addr[2884] = 382;
        test_data[2884] = 33'd8361796239;
        test_addr[2885] = 383;
        test_data[2885] = 33'd6335079144;
        test_addr[2886] = 384;
        test_data[2886] = 33'd6969592656;
        test_addr[2887] = 385;
        test_data[2887] = 33'd817202464;
        test_addr[2888] = 386;
        test_data[2888] = 33'd3041406532;
        test_addr[2889] = 387;
        test_data[2889] = 33'd1591272145;
        test_addr[2890] = 388;
        test_data[2890] = 33'd4926402922;
        test_addr[2891] = 389;
        test_data[2891] = 33'd3497432784;
        test_addr[2892] = 390;
        test_data[2892] = 33'd2543760664;
        test_addr[2893] = 8;
        test_data[2893] = 33'd3378399337;
        test_addr[2894] = 9;
        test_data[2894] = 33'd1114041214;
        test_addr[2895] = 10;
        test_data[2895] = 33'd8228532721;
        test_addr[2896] = 11;
        test_data[2896] = 33'd874847442;
        test_addr[2897] = 12;
        test_data[2897] = 33'd5729417136;
        test_addr[2898] = 13;
        test_data[2898] = 33'd2440374455;
        test_addr[2899] = 14;
        test_data[2899] = 33'd7725903567;
        test_addr[2900] = 15;
        test_data[2900] = 33'd3854493493;
        test_addr[2901] = 391;
        test_data[2901] = 33'd189757725;
        test_addr[2902] = 392;
        test_data[2902] = 33'd6383939894;
        test_addr[2903] = 393;
        test_data[2903] = 33'd8553094591;
        test_addr[2904] = 394;
        test_data[2904] = 33'd4845477181;
        test_addr[2905] = 395;
        test_data[2905] = 33'd1735085298;
        test_addr[2906] = 396;
        test_data[2906] = 33'd5758080572;
        test_addr[2907] = 397;
        test_data[2907] = 33'd4140998441;
        test_addr[2908] = 398;
        test_data[2908] = 33'd3505084960;
        test_addr[2909] = 399;
        test_data[2909] = 33'd5856656725;
        test_addr[2910] = 400;
        test_data[2910] = 33'd8462755297;
        test_addr[2911] = 853;
        test_data[2911] = 33'd1067052146;
        test_addr[2912] = 854;
        test_data[2912] = 33'd5159156605;
        test_addr[2913] = 855;
        test_data[2913] = 33'd1604534845;
        test_addr[2914] = 856;
        test_data[2914] = 33'd821537468;
        test_addr[2915] = 857;
        test_data[2915] = 33'd179268970;
        test_addr[2916] = 858;
        test_data[2916] = 33'd724552190;
        test_addr[2917] = 859;
        test_data[2917] = 33'd6222611576;
        test_addr[2918] = 860;
        test_data[2918] = 33'd9740189;
        test_addr[2919] = 861;
        test_data[2919] = 33'd4244904036;
        test_addr[2920] = 862;
        test_data[2920] = 33'd4180459732;
        test_addr[2921] = 863;
        test_data[2921] = 33'd3181973309;
        test_addr[2922] = 864;
        test_data[2922] = 33'd4122567500;
        test_addr[2923] = 865;
        test_data[2923] = 33'd2442557656;
        test_addr[2924] = 866;
        test_data[2924] = 33'd636310232;
        test_addr[2925] = 867;
        test_data[2925] = 33'd6977750975;
        test_addr[2926] = 401;
        test_data[2926] = 33'd427139017;
        test_addr[2927] = 402;
        test_data[2927] = 33'd1203385049;
        test_addr[2928] = 403;
        test_data[2928] = 33'd534753598;
        test_addr[2929] = 404;
        test_data[2929] = 33'd128960265;
        test_addr[2930] = 520;
        test_data[2930] = 33'd5852278765;
        test_addr[2931] = 521;
        test_data[2931] = 33'd4960232593;
        test_addr[2932] = 522;
        test_data[2932] = 33'd3048636483;
        test_addr[2933] = 523;
        test_data[2933] = 33'd1382851467;
        test_addr[2934] = 524;
        test_data[2934] = 33'd8038907190;
        test_addr[2935] = 525;
        test_data[2935] = 33'd2281015751;
        test_addr[2936] = 526;
        test_data[2936] = 33'd5969965825;
        test_addr[2937] = 527;
        test_data[2937] = 33'd3884199812;
        test_addr[2938] = 405;
        test_data[2938] = 33'd4388752602;
        test_addr[2939] = 406;
        test_data[2939] = 33'd4270269366;
        test_addr[2940] = 407;
        test_data[2940] = 33'd3650981421;
        test_addr[2941] = 408;
        test_data[2941] = 33'd1991242564;
        test_addr[2942] = 409;
        test_data[2942] = 33'd881702054;
        test_addr[2943] = 363;
        test_data[2943] = 33'd2723076636;
        test_addr[2944] = 364;
        test_data[2944] = 33'd1714130166;
        test_addr[2945] = 365;
        test_data[2945] = 33'd6996148361;
        test_addr[2946] = 366;
        test_data[2946] = 33'd1589586476;
        test_addr[2947] = 367;
        test_data[2947] = 33'd3426483264;
        test_addr[2948] = 410;
        test_data[2948] = 33'd3442998655;
        test_addr[2949] = 411;
        test_data[2949] = 33'd1375207748;
        test_addr[2950] = 412;
        test_data[2950] = 33'd5360105389;
        test_addr[2951] = 413;
        test_data[2951] = 33'd6660651092;
        test_addr[2952] = 414;
        test_data[2952] = 33'd2622463751;
        test_addr[2953] = 415;
        test_data[2953] = 33'd2483981373;
        test_addr[2954] = 416;
        test_data[2954] = 33'd3762483973;
        test_addr[2955] = 417;
        test_data[2955] = 33'd857483597;
        test_addr[2956] = 418;
        test_data[2956] = 33'd3304050455;
        test_addr[2957] = 419;
        test_data[2957] = 33'd8558011129;
        test_addr[2958] = 420;
        test_data[2958] = 33'd2008269494;
        test_addr[2959] = 421;
        test_data[2959] = 33'd3124744987;
        test_addr[2960] = 422;
        test_data[2960] = 33'd5526307217;
        test_addr[2961] = 423;
        test_data[2961] = 33'd3101606753;
        test_addr[2962] = 424;
        test_data[2962] = 33'd4107482093;
        test_addr[2963] = 425;
        test_data[2963] = 33'd2446718652;
        test_addr[2964] = 999;
        test_data[2964] = 33'd5525547260;
        test_addr[2965] = 1000;
        test_data[2965] = 33'd4512195154;
        test_addr[2966] = 1001;
        test_data[2966] = 33'd1757685921;
        test_addr[2967] = 1002;
        test_data[2967] = 33'd1476013580;
        test_addr[2968] = 1003;
        test_data[2968] = 33'd6928504097;
        test_addr[2969] = 1004;
        test_data[2969] = 33'd3198229176;
        test_addr[2970] = 1005;
        test_data[2970] = 33'd2395804748;
        test_addr[2971] = 1006;
        test_data[2971] = 33'd4558578965;
        test_addr[2972] = 1007;
        test_data[2972] = 33'd4059948122;
        test_addr[2973] = 1008;
        test_data[2973] = 33'd7341823353;
        test_addr[2974] = 1009;
        test_data[2974] = 33'd2905712961;
        test_addr[2975] = 1010;
        test_data[2975] = 33'd7083158790;
        test_addr[2976] = 1011;
        test_data[2976] = 33'd6638230579;
        test_addr[2977] = 1012;
        test_data[2977] = 33'd4866929644;
        test_addr[2978] = 1013;
        test_data[2978] = 33'd1050220471;
        test_addr[2979] = 1014;
        test_data[2979] = 33'd460798996;
        test_addr[2980] = 1015;
        test_data[2980] = 33'd6525946098;
        test_addr[2981] = 1016;
        test_data[2981] = 33'd3061783049;
        test_addr[2982] = 1017;
        test_data[2982] = 33'd293708126;
        test_addr[2983] = 1018;
        test_data[2983] = 33'd7412945313;
        test_addr[2984] = 1019;
        test_data[2984] = 33'd1738985240;
        test_addr[2985] = 1020;
        test_data[2985] = 33'd1804380535;
        test_addr[2986] = 1021;
        test_data[2986] = 33'd1888120797;
        test_addr[2987] = 1022;
        test_data[2987] = 33'd1248002737;
        test_addr[2988] = 1023;
        test_data[2988] = 33'd3674196659;
        test_addr[2989] = 0;
        test_data[2989] = 33'd8215530205;
        test_addr[2990] = 1;
        test_data[2990] = 33'd1869574933;
        test_addr[2991] = 2;
        test_data[2991] = 33'd728813621;
        test_addr[2992] = 3;
        test_data[2992] = 33'd7625901397;
        test_addr[2993] = 4;
        test_data[2993] = 33'd4417781632;
        test_addr[2994] = 5;
        test_data[2994] = 33'd485978242;
        test_addr[2995] = 6;
        test_data[2995] = 33'd4875743580;
        test_addr[2996] = 7;
        test_data[2996] = 33'd4602426284;
        test_addr[2997] = 8;
        test_data[2997] = 33'd5408630530;
        test_addr[2998] = 9;
        test_data[2998] = 33'd1114041214;
        test_addr[2999] = 426;
        test_data[2999] = 33'd3096364448;

    end
endmodule
